magic
tech sky130A
magscale 1 2
timestamp 1725190886
<< nwell >>
rect 24100 -4757 24530 -4756
rect 19257 -5355 19445 -5352
rect 20362 -5355 20676 -5352
rect 18919 -5358 20676 -5355
rect 18919 -7120 20883 -5358
rect 24100 -6921 24702 -4757
rect 26205 -6494 26499 -4753
rect 26188 -6918 26499 -6494
rect 19257 -7127 20883 -7120
<< pwell >>
rect 23148 -7850 23290 -7798
rect 23884 -7845 23954 -7746
rect 24974 -7845 25044 -7739
rect 25638 -7873 25708 -7823
rect 25804 -7856 26040 -7832
rect 25947 -7995 26008 -7856
rect 23071 -8122 23136 -8091
rect 23140 -8878 23190 -8621
rect 25947 -8685 26031 -7995
rect 25947 -8874 26008 -8685
rect 24216 -8978 24286 -8877
rect 25306 -8909 25376 -8877
rect 25306 -8953 25420 -8909
rect 25804 -8910 26040 -8874
rect 25306 -8978 25376 -8953
rect 26048 -9258 26072 -9227
rect 23058 -9708 23337 -9297
rect 25668 -9360 25669 -9260
rect 25784 -9394 26072 -9258
rect 23060 -9808 23127 -9708
rect 26048 -9947 26072 -9394
rect 23105 -10359 23326 -9964
rect 25782 -10512 26042 -10332
<< nbase >>
rect 29575 -9292 29614 -9291
<< pdiff >>
rect 29575 -9292 29614 -9291
<< psubdiff >>
rect 16171 -3802 16195 -3600
rect 33602 -3802 33626 -3600
rect 16200 -4004 16402 -3980
rect 33402 -4202 33606 -4178
rect 16900 -7475 17099 -7399
rect 16900 -8923 16943 -7475
rect 17049 -8923 17099 -7475
rect 16900 -9000 17099 -8923
rect 22599 -7469 22798 -7393
rect 22599 -8917 22642 -7469
rect 22748 -8917 22798 -7469
rect 22599 -8992 22798 -8917
rect 22726 -8996 22798 -8992
rect 19198 -9426 19404 -9399
rect 19198 -9787 19258 -9426
rect 19323 -9787 19404 -9426
rect 19198 -9800 19404 -9787
rect 20500 -9421 20705 -9394
rect 20500 -9782 20559 -9421
rect 20624 -9782 20705 -9421
rect 20500 -9795 20705 -9782
rect 33402 -12426 33606 -12402
rect 16200 -12624 16402 -12600
rect 16172 -12997 16196 -12799
rect 33598 -12997 33622 -12799
<< nsubdiff >>
rect 24300 -4967 24403 -4901
rect 19067 -5457 19216 -5403
rect 19067 -6902 19097 -5457
rect 19184 -6902 19216 -5457
rect 19067 -7004 19216 -6902
rect 20500 -5457 20649 -5398
rect 20500 -6902 20528 -5457
rect 20615 -6902 20649 -5457
rect 24300 -6747 24329 -4967
rect 24372 -6747 24403 -4967
rect 24300 -6802 24403 -6747
rect 26305 -4967 26408 -4901
rect 26305 -6747 26334 -4967
rect 26377 -6747 26408 -4967
rect 26305 -6802 26408 -6747
rect 20500 -6999 20649 -6902
<< psubdiffcont >>
rect 16195 -3802 33602 -3600
rect 16200 -12600 16402 -4004
rect 16943 -8923 17049 -7475
rect 22642 -8917 22748 -7469
rect 19258 -9787 19323 -9426
rect 20559 -9782 20624 -9421
rect 33402 -12402 33606 -4202
rect 16196 -12997 33598 -12799
<< nsubdiffcont >>
rect 19097 -6902 19184 -5457
rect 20528 -6902 20615 -5457
rect 24329 -6747 24372 -4967
rect 26334 -6747 26377 -4967
<< locali >>
rect 16179 -3802 16195 -3600
rect 33602 -3802 33618 -3600
rect 16202 -3988 16402 -3802
rect 16200 -4004 16402 -3988
rect 33400 -4100 33602 -3802
rect 33400 -4174 33606 -4100
rect 33402 -4202 33606 -4174
rect 26630 -4488 33006 -4471
rect 26630 -4707 33070 -4488
rect 19084 -5430 19197 -5429
rect 20518 -5434 20631 -5433
rect 19197 -5969 19198 -5467
rect 19084 -6902 19097 -6182
rect 19184 -6902 19197 -6182
rect 19084 -6954 19197 -6902
rect 20518 -6052 20521 -5434
rect 20518 -6902 20528 -6052
rect 20615 -6902 20631 -6052
rect 24317 -6221 24329 -5200
rect 24372 -6221 24384 -5200
rect 24317 -6720 24319 -6221
rect 26322 -6225 26334 -5200
rect 26377 -6225 26389 -5200
rect 26631 -5996 33071 -5523
rect 24317 -6747 24329 -6720
rect 24372 -6747 24384 -6720
rect 24317 -6784 24384 -6747
rect 26322 -6747 26334 -6724
rect 26377 -6747 26389 -6724
rect 26322 -6784 26389 -6747
rect 20518 -6958 20631 -6902
rect 26630 -7284 33073 -6813
rect 16929 -7475 17070 -7444
rect 16929 -8923 16943 -7475
rect 17049 -8923 17070 -7475
rect 22628 -7469 22769 -7438
rect 16929 -8926 16960 -8923
rect 17029 -8926 17070 -8923
rect 16929 -8973 17070 -8926
rect 22628 -8917 22642 -7469
rect 22748 -8917 22769 -7469
rect 26627 -8572 33072 -8099
rect 22628 -8967 22769 -8917
rect 29575 -9292 29614 -9291
rect 19242 -9426 19348 -9401
rect 19242 -9787 19258 -9426
rect 19323 -9787 19348 -9426
rect 19242 -9804 19348 -9787
rect 20543 -9421 20649 -9396
rect 20543 -9782 20559 -9421
rect 20624 -9782 20649 -9421
rect 20543 -9799 20649 -9782
rect 26625 -9792 33073 -9388
rect 32669 -9861 33073 -9792
rect 26006 -10357 26043 -10331
rect 32660 -10732 33072 -10676
rect 26626 -11146 33073 -10732
rect 26635 -12182 33065 -11964
rect 26635 -12199 33006 -12182
rect 16200 -12616 16402 -12600
rect 16202 -12799 16402 -12616
rect 33400 -12418 33606 -12402
rect 33400 -12799 33598 -12418
rect 16180 -12997 16196 -12799
rect 33598 -12997 33614 -12799
rect 16202 -13000 16402 -12997
<< viali >>
rect 19083 -5457 19197 -5430
rect 19083 -6182 19097 -5457
rect 19097 -6182 19184 -5457
rect 19184 -6182 19197 -5457
rect 20521 -5457 20634 -5434
rect 20521 -6052 20528 -5457
rect 20528 -6052 20615 -5457
rect 20615 -6052 20634 -5457
rect 21440 -6577 21498 -4880
rect 24316 -4967 24386 -4932
rect 24316 -5200 24329 -4967
rect 24329 -5200 24372 -4967
rect 24372 -5200 24386 -4967
rect 26320 -4967 26390 -4898
rect 26320 -5166 26334 -4967
rect 26334 -5166 26377 -4967
rect 26377 -5166 26390 -4967
rect 24319 -6720 24329 -6221
rect 24329 -6720 24372 -6221
rect 24372 -6720 24387 -6221
rect 26321 -6724 26334 -6225
rect 26334 -6724 26377 -6225
rect 26377 -6724 26389 -6225
rect 16204 -7774 16402 -7506
rect 16402 -7774 16468 -7506
rect 16960 -8923 17029 -7506
rect 18012 -7800 18048 -7512
rect 21674 -7802 21718 -7550
rect 16960 -8926 17029 -8923
rect 22655 -8909 22724 -7489
rect 23717 -7749 23789 -7715
rect 23087 -8065 23128 -7834
rect 25969 -8099 26004 -7845
rect 23089 -8845 23130 -8614
rect 25969 -8876 26004 -8622
rect 23385 -9007 23456 -8973
rect 19258 -9557 19323 -9426
rect 19258 -9787 19323 -9650
rect 20559 -9552 20624 -9421
rect 20559 -9782 20624 -9645
rect 23060 -9698 23097 -9305
rect 26005 -9700 26042 -9307
rect 23068 -10358 23105 -9965
rect 26006 -10331 26043 -9964
rect 23038 -12985 23152 -12871
rect 25954 -12987 26068 -12873
<< metal1 >>
rect 22344 -4257 26216 -4255
rect 22344 -4385 26158 -4257
rect 22344 -4388 22550 -4385
rect 26152 -4388 26158 -4385
rect 26289 -4388 26295 -4257
rect 22344 -4496 22549 -4388
rect 21407 -4880 21610 -4745
rect 22343 -4854 22549 -4496
rect 24195 -4502 25934 -4500
rect 24068 -4631 24074 -4502
rect 24203 -4596 25934 -4502
rect 24203 -4631 25935 -4596
rect 24195 -4696 25935 -4631
rect 24201 -4700 25935 -4696
rect 24768 -4755 25935 -4700
rect 24323 -4815 24694 -4755
rect 24753 -4815 25959 -4755
rect 26018 -4815 26386 -4755
rect 19640 -5363 20104 -5357
rect 19077 -5430 19203 -5418
rect 19640 -5426 19700 -5363
rect 19073 -5536 19083 -5430
rect 19070 -5856 19083 -5536
rect 19073 -6182 19083 -5856
rect 19197 -5536 19207 -5430
rect 19694 -5465 19700 -5426
rect 19802 -5426 20104 -5363
rect 19802 -5465 19808 -5426
rect 20515 -5434 20640 -5422
rect 20511 -5536 20521 -5434
rect 19197 -5856 20521 -5536
rect 19197 -6182 19207 -5856
rect 20511 -6052 20521 -5856
rect 20634 -6052 20644 -5434
rect 20515 -6064 20640 -6052
rect 19077 -6194 19203 -6182
rect 19538 -6571 19667 -6530
rect 19538 -6673 19563 -6571
rect 19665 -6673 19667 -6571
rect 18964 -7038 19093 -7037
rect 19538 -7038 19667 -6673
rect 18964 -7167 19667 -7038
rect 20073 -7042 20202 -6534
rect 21407 -6573 21440 -4880
rect 21406 -6577 21440 -6573
rect 21498 -6573 21610 -4880
rect 22104 -6570 23116 -4854
rect 24323 -4879 24383 -4815
rect 26326 -4878 26386 -4815
rect 26292 -4879 26412 -4878
rect 24299 -4880 26412 -4879
rect 24298 -4898 26412 -4880
rect 24298 -4932 26320 -4898
rect 21498 -6577 21671 -6573
rect 21406 -6912 21671 -6577
rect 23614 -6775 23668 -4961
rect 24298 -5200 24316 -4932
rect 24386 -5166 26320 -4932
rect 26390 -5166 26412 -4898
rect 24386 -5200 26412 -5166
rect 24298 -5204 26412 -5200
rect 24298 -5206 24412 -5204
rect 26288 -5206 26412 -5204
rect 24298 -5208 24402 -5206
rect 24310 -5212 24392 -5208
rect 25775 -5976 26035 -5975
rect 26158 -5976 26288 -5970
rect 25775 -6106 26158 -5976
rect 24313 -6220 24393 -6209
rect 24308 -6720 24318 -6220
rect 24388 -6720 24590 -6220
rect 24313 -6732 24393 -6720
rect 22666 -6829 23668 -6775
rect 21406 -6913 21764 -6912
rect 21406 -7040 22468 -6913
rect 22595 -7040 22601 -6913
rect 20752 -7041 21086 -7040
rect 20647 -7042 21086 -7041
rect 20073 -7070 21086 -7042
rect 21406 -7070 22249 -7040
rect 20073 -7163 22249 -7070
rect 16954 -7495 17035 -7494
rect 16343 -7500 17106 -7495
rect 16192 -7502 17309 -7500
rect 16192 -7506 17317 -7502
rect 16192 -7774 16204 -7506
rect 16468 -7774 16960 -7506
rect 16192 -7780 16960 -7774
rect 16343 -7789 16960 -7780
rect 16946 -7801 16960 -7789
rect 16954 -8926 16960 -7801
rect 17029 -7513 17317 -7506
rect 18006 -7512 18054 -7500
rect 18006 -7513 18012 -7512
rect 17029 -7800 18012 -7513
rect 18048 -7513 18054 -7512
rect 18048 -7800 18080 -7513
rect 17029 -7801 18080 -7800
rect 17029 -8926 17035 -7801
rect 17188 -7803 17317 -7801
rect 18006 -7812 18054 -7801
rect 18964 -7888 19093 -7167
rect 20073 -7171 21086 -7163
rect 21630 -7164 22249 -7163
rect 20647 -7172 21086 -7171
rect 20647 -7892 20776 -7172
rect 22666 -7469 22720 -6829
rect 24816 -7158 24944 -6218
rect 22830 -7277 24944 -7158
rect 22666 -7477 22724 -7469
rect 22649 -7489 22730 -7477
rect 21620 -7502 22404 -7500
rect 22649 -7502 22655 -7489
rect 21620 -7550 22655 -7502
rect 21620 -7802 21674 -7550
rect 21718 -7802 22655 -7550
rect 21668 -7814 21724 -7802
rect 22403 -7803 22655 -7802
rect 22649 -8099 22655 -7803
rect 22636 -8340 22655 -8099
rect 19829 -8446 19839 -8445
rect 18126 -8701 19839 -8446
rect 19905 -8446 19915 -8445
rect 19905 -8447 21608 -8446
rect 19905 -8701 21609 -8447
rect 22649 -8589 22655 -8340
rect 21584 -8710 21609 -8701
rect 22626 -8875 22655 -8589
rect 22630 -8909 22655 -8875
rect 22724 -8099 22730 -7489
rect 22830 -7569 22964 -7277
rect 24904 -7278 24944 -7277
rect 25146 -7183 25255 -6220
rect 25146 -7558 25255 -7292
rect 25454 -7387 25563 -6215
rect 25775 -7089 25893 -6106
rect 26158 -6112 26288 -6106
rect 26315 -6224 26395 -6213
rect 26132 -6723 26320 -6224
rect 26392 -6723 26402 -6224
rect 26132 -6724 26321 -6723
rect 26389 -6724 26402 -6723
rect 26315 -6736 26395 -6724
rect 25775 -7207 26289 -7089
rect 25454 -7502 25563 -7496
rect 24520 -7568 25708 -7558
rect 22823 -7703 22829 -7569
rect 22963 -7703 22969 -7569
rect 24519 -7620 24525 -7568
rect 24577 -7620 25708 -7568
rect 24520 -7628 25708 -7620
rect 23705 -7715 23801 -7709
rect 23705 -7749 23717 -7715
rect 23789 -7749 23801 -7715
rect 23705 -7755 23801 -7749
rect 23148 -7799 23290 -7798
rect 23053 -7800 23290 -7799
rect 23033 -7834 23290 -7800
rect 23033 -8065 23087 -7834
rect 23128 -8065 23290 -7834
rect 22724 -8340 22770 -8099
rect 23033 -8100 23290 -8065
rect 23386 -7845 23456 -7844
rect 23386 -8001 23622 -7845
rect 22724 -8589 22730 -8340
rect 23033 -8469 23149 -8100
rect 23386 -8277 23456 -8001
rect 23552 -8278 23622 -8001
rect 23717 -8277 23789 -7755
rect 23884 -7809 24878 -7739
rect 23884 -8278 23954 -7809
rect 24049 -8001 24286 -7845
rect 24049 -8278 24119 -8001
rect 24216 -8278 24286 -8001
rect 24528 -8187 24577 -7880
rect 24519 -8239 24525 -8187
rect 24577 -8239 24583 -8187
rect 24528 -8246 24577 -8239
rect 24808 -8278 24878 -7809
rect 24974 -7809 25542 -7739
rect 24974 -8278 25044 -7809
rect 25140 -8001 25376 -7845
rect 25140 -8278 25210 -8001
rect 25306 -8278 25376 -8001
rect 25472 -8278 25542 -7809
rect 25638 -8277 25708 -7628
rect 25804 -7845 26040 -7832
rect 25804 -8099 25969 -7845
rect 26004 -8099 26040 -7845
rect 25804 -8100 26040 -8099
rect 24511 -8422 24517 -8417
rect 23032 -8567 23149 -8469
rect 23032 -8588 23150 -8567
rect 23032 -8589 23290 -8588
rect 22724 -8614 23290 -8589
rect 22724 -8845 23089 -8614
rect 23130 -8845 23290 -8614
rect 22724 -8875 23290 -8845
rect 22724 -8909 22792 -8875
rect 22630 -8918 22792 -8909
rect 23032 -8877 23290 -8875
rect 23032 -8878 23190 -8877
rect 16954 -8938 17035 -8926
rect 16964 -8974 17028 -8938
rect 19694 -8992 19704 -8960
rect 18181 -9048 19704 -8992
rect 19800 -9048 19810 -8960
rect 19990 -8992 20000 -8960
rect 19931 -9048 20000 -8992
rect 20100 -8992 20110 -8960
rect 20100 -9048 21555 -8992
rect 19835 -9247 19841 -9187
rect 19901 -9247 19907 -9187
rect 19252 -9421 19329 -9414
rect 19252 -9426 19578 -9421
rect 19252 -9557 19258 -9426
rect 19323 -9557 19578 -9426
rect 19252 -9558 19578 -9557
rect 19252 -9569 19329 -9558
rect 19841 -9561 19901 -9247
rect 20155 -9309 22829 -9175
rect 22963 -9309 22969 -9175
rect 23032 -9297 23149 -8878
rect 23385 -8967 23456 -8501
rect 23552 -8906 23622 -8443
rect 23884 -8721 23954 -8443
rect 23718 -8877 23954 -8721
rect 24049 -8906 24119 -8443
rect 23373 -8973 23468 -8967
rect 23373 -9007 23385 -8973
rect 23456 -9007 23468 -8973
rect 23552 -8976 24119 -8906
rect 24216 -8908 24286 -8443
rect 24509 -8473 24517 -8422
rect 24573 -8422 24579 -8417
rect 24573 -8473 24584 -8422
rect 24509 -8830 24584 -8473
rect 24808 -8721 24878 -8436
rect 24974 -8721 25044 -8436
rect 24808 -8877 25044 -8721
rect 24808 -8878 24878 -8877
rect 25140 -8908 25210 -8436
rect 24216 -8978 25210 -8908
rect 25306 -8903 25376 -8447
rect 25472 -8721 25542 -8436
rect 25947 -8622 26040 -8100
rect 25472 -8877 25708 -8721
rect 25804 -8876 25969 -8622
rect 26004 -8876 26040 -8622
rect 25358 -8955 25376 -8903
rect 25804 -8910 26040 -8876
rect 25306 -8972 25376 -8955
rect 23373 -9013 23468 -9007
rect 26171 -9060 26289 -7207
rect 25551 -9131 26289 -9060
rect 25549 -9178 26289 -9131
rect 26925 -7285 32772 -4768
rect 26925 -8098 29439 -7285
rect 29528 -7600 30172 -7382
rect 29528 -7802 29809 -7600
rect 30011 -7802 30172 -7600
rect 29528 -8006 30172 -7802
rect 30255 -8098 32772 -7285
rect 26925 -8749 32772 -8098
rect 26925 -8799 29547 -8749
rect 29578 -8799 32772 -8749
rect 26925 -9000 32772 -8799
rect 25549 -9217 25916 -9178
rect 26925 -9200 29807 -9000
rect 30007 -9200 32772 -9000
rect 23032 -9305 23337 -9297
rect 19252 -9650 19348 -9638
rect 19227 -9787 19258 -9650
rect 19323 -9787 20057 -9650
rect 20155 -9747 20217 -9309
rect 20553 -9416 20630 -9409
rect 20553 -9421 20649 -9416
rect 20553 -9552 20559 -9421
rect 20624 -9552 20649 -9421
rect 20553 -9553 20649 -9552
rect 20553 -9564 20630 -9553
rect 19252 -9793 19348 -9787
rect 19252 -9799 19341 -9793
rect 19684 -9794 19774 -9787
rect 19276 -9836 19341 -9799
rect 20095 -9809 20217 -9747
rect 20315 -9645 20651 -9632
rect 20315 -9782 20559 -9645
rect 20624 -9653 20651 -9645
rect 20624 -9782 20652 -9653
rect 20315 -9797 20652 -9782
rect 23032 -9698 23060 -9305
rect 23097 -9310 23337 -9305
rect 23445 -9310 23564 -9297
rect 23097 -9698 23564 -9310
rect 23032 -9707 23564 -9698
rect 23032 -9708 23337 -9707
rect 20315 -9808 20651 -9797
rect 19276 -9899 19687 -9836
rect 20095 -9841 20157 -9809
rect 20519 -9837 20651 -9808
rect 19741 -9899 20158 -9841
rect 20211 -9893 20651 -9837
rect 19399 -10134 19510 -9899
rect 20216 -10134 20327 -9893
rect 19399 -10245 20327 -10134
rect 23032 -9964 23149 -9708
rect 23445 -9725 23564 -9707
rect 23677 -9310 23796 -9299
rect 23912 -9310 24031 -9297
rect 23677 -9707 24031 -9310
rect 23677 -9725 23796 -9707
rect 23912 -9725 24031 -9707
rect 24147 -9313 24266 -9297
rect 24381 -9313 24500 -9298
rect 24147 -9710 24500 -9313
rect 24147 -9725 24266 -9710
rect 24381 -9725 24500 -9710
rect 24614 -9308 24733 -9298
rect 24848 -9308 24967 -9297
rect 24614 -9705 24967 -9308
rect 24614 -9725 24733 -9705
rect 24848 -9725 24967 -9705
rect 25083 -9311 25202 -9298
rect 25316 -9311 25435 -9298
rect 25083 -9708 25435 -9311
rect 25549 -9582 25669 -9217
rect 25784 -9261 26064 -9258
rect 25784 -9307 26074 -9261
rect 25784 -9394 26005 -9307
rect 25083 -9725 25202 -9708
rect 25316 -9725 25435 -9708
rect 25550 -9719 25669 -9582
rect 25790 -9700 26005 -9394
rect 26042 -9700 26074 -9307
rect 25790 -9705 26074 -9700
rect 23445 -9961 23564 -9945
rect 23677 -9961 23796 -9942
rect 23032 -9965 23326 -9964
rect 23032 -10358 23068 -9965
rect 23105 -10358 23326 -9965
rect 23032 -10359 23326 -10358
rect 23445 -10358 23796 -9961
rect 23032 -12871 23158 -10359
rect 23445 -10370 23564 -10358
rect 23677 -10372 23796 -10358
rect 23912 -9961 24031 -9942
rect 24147 -9961 24266 -9942
rect 23912 -10358 24266 -9961
rect 23912 -10370 24031 -10358
rect 24147 -10370 24266 -10358
rect 24381 -9961 24500 -9942
rect 24614 -9961 24733 -9942
rect 24381 -10358 24733 -9961
rect 24381 -10371 24500 -10358
rect 24614 -10371 24733 -10358
rect 24848 -9961 24967 -9942
rect 25083 -9961 25202 -9942
rect 24848 -10358 25202 -9961
rect 24848 -10370 24967 -10358
rect 25083 -10371 25202 -10358
rect 25316 -9963 25435 -9942
rect 25550 -9963 25669 -9945
rect 25981 -9963 26074 -9705
rect 25316 -10360 25669 -9963
rect 25789 -9964 26074 -9963
rect 25789 -10331 26006 -9964
rect 26043 -10331 26074 -9964
rect 25789 -10332 26074 -10331
rect 25316 -10371 25435 -10360
rect 25550 -10372 25669 -10360
rect 25782 -10512 26074 -10332
rect 23032 -12985 23038 -12871
rect 23152 -12985 23158 -12871
rect 23032 -12997 23158 -12985
rect 25948 -12873 26074 -10512
rect 26925 -11902 32772 -9200
rect 25948 -12987 25954 -12873
rect 26068 -12987 26074 -12873
rect 25948 -12999 26074 -12987
<< via1 >>
rect 26158 -4388 26289 -4257
rect 24074 -4631 24203 -4502
rect 19083 -6182 19197 -5430
rect 19700 -5465 19802 -5363
rect 20521 -6052 20634 -5434
rect 19563 -6673 19665 -6571
rect 24316 -5200 24386 -4932
rect 26320 -5166 26390 -4898
rect 26158 -6106 26288 -5976
rect 24318 -6221 24388 -6220
rect 24318 -6720 24319 -6221
rect 24319 -6720 24387 -6221
rect 24387 -6720 24388 -6221
rect 22468 -7040 22595 -6913
rect 19839 -8701 19905 -8445
rect 25146 -7292 25255 -7183
rect 26320 -6225 26392 -6224
rect 26320 -6723 26321 -6225
rect 26321 -6723 26389 -6225
rect 26389 -6723 26392 -6225
rect 25454 -7496 25563 -7387
rect 22829 -7703 22963 -7569
rect 24525 -7620 24577 -7568
rect 24525 -8239 24577 -8187
rect 19704 -9048 19800 -8960
rect 20000 -9048 20100 -8960
rect 19841 -9247 19901 -9187
rect 22829 -9309 22963 -9175
rect 24517 -8473 24573 -8417
rect 25306 -8955 25358 -8903
rect 29809 -7802 30011 -7600
rect 29807 -9200 30007 -9000
<< metal2 >>
rect 26158 -4257 26289 -4251
rect 24074 -4502 24203 -4496
rect 19700 -5363 19802 -5357
rect 19083 -5430 19197 -5420
rect 19083 -6192 19197 -6182
rect 19700 -6571 19802 -5465
rect 20521 -5434 20634 -5424
rect 20521 -6062 20634 -6052
rect 19557 -6673 19563 -6571
rect 19665 -6673 19802 -6571
rect 22468 -6910 22595 -6907
rect 24074 -6910 24203 -4631
rect 24316 -4932 24386 -4922
rect 24316 -5210 24386 -5200
rect 26158 -5976 26289 -4388
rect 26320 -4898 26390 -4888
rect 26320 -5176 26390 -5166
rect 26152 -6106 26158 -5976
rect 26288 -6106 26294 -5976
rect 24318 -6220 24388 -6210
rect 24318 -6730 24388 -6720
rect 26320 -6224 26392 -6214
rect 26320 -6733 26392 -6723
rect 22468 -6913 24203 -6910
rect 22595 -7040 24203 -6913
rect 22468 -7046 22595 -7040
rect 25140 -7199 25146 -7183
rect 19704 -7292 25146 -7199
rect 25255 -7292 25261 -7183
rect 19704 -7299 25261 -7292
rect 19704 -8960 19804 -7299
rect 25448 -7397 25454 -7387
rect 20001 -7496 25454 -7397
rect 25563 -7397 25569 -7387
rect 26402 -7397 26604 -7394
rect 25563 -7496 26604 -7397
rect 20001 -7497 26604 -7496
rect 19839 -8445 19905 -8435
rect 19839 -8711 19905 -8701
rect 19840 -8950 19902 -8711
rect 20001 -8950 20101 -7497
rect 19800 -9040 19804 -8960
rect 19704 -9058 19800 -9048
rect 19841 -9187 19901 -8950
rect 20000 -8960 20101 -8950
rect 20100 -9043 20101 -8960
rect 22829 -7569 22963 -7563
rect 22829 -8073 22963 -7703
rect 24514 -7568 24599 -7555
rect 24514 -7620 24525 -7568
rect 24577 -7620 24599 -7568
rect 22829 -8451 22964 -8073
rect 24514 -8187 24599 -7620
rect 24514 -8239 24525 -8187
rect 24577 -8239 24599 -8187
rect 24514 -8257 24599 -8239
rect 24517 -8417 24573 -8411
rect 20000 -9058 20100 -9048
rect 19841 -9253 19901 -9247
rect 22829 -9175 22963 -8451
rect 24517 -9006 24573 -8473
rect 25300 -8955 25306 -8903
rect 25358 -8905 25364 -8903
rect 25461 -8905 25555 -7497
rect 26402 -7600 26604 -7497
rect 26402 -7802 29809 -7600
rect 30011 -7802 30017 -7600
rect 25358 -8953 25555 -8905
rect 25358 -8955 25364 -8953
rect 25400 -8955 25555 -8953
rect 26400 -9000 26799 -8999
rect 26400 -9006 29807 -9000
rect 24517 -9196 29807 -9006
rect 26400 -9200 29807 -9196
rect 30007 -9200 30013 -9000
rect 22829 -9315 22963 -9309
<< via2 >>
rect 19083 -6182 19197 -5430
rect 20521 -6052 20634 -5434
rect 24316 -5200 24386 -4932
rect 26320 -5166 26390 -4898
rect 24318 -6720 24388 -6220
rect 26320 -6723 26392 -6224
<< metal3 >>
rect 20616 -4526 26396 -4525
rect 19095 -4704 26396 -4526
rect 19095 -4882 20636 -4704
rect 19101 -5425 19215 -4882
rect 19073 -5430 19215 -5425
rect 20532 -5429 20636 -4882
rect 24312 -4927 24384 -4704
rect 26320 -4893 26392 -4704
rect 26310 -4898 26400 -4893
rect 24306 -4932 24396 -4927
rect 24306 -5200 24316 -4932
rect 24386 -5200 24396 -4932
rect 26310 -5166 26320 -4898
rect 26390 -5166 26400 -4898
rect 26310 -5171 26400 -5166
rect 24306 -5205 24396 -5200
rect 19073 -6182 19083 -5430
rect 19197 -5494 19215 -5430
rect 20511 -5434 20644 -5429
rect 19197 -6182 19207 -5494
rect 20511 -6052 20521 -5434
rect 20634 -6052 20644 -5434
rect 20511 -6057 20644 -6052
rect 19073 -6187 19207 -6182
rect 24312 -6215 24384 -5205
rect 24308 -6220 24398 -6215
rect 26320 -6219 26392 -5171
rect 24308 -6720 24318 -6220
rect 24388 -6720 24398 -6220
rect 24308 -6725 24398 -6720
rect 26310 -6224 26402 -6219
rect 26310 -6723 26320 -6224
rect 26392 -6723 26402 -6224
rect 24312 -6729 24384 -6725
rect 26310 -6728 26402 -6723
rect 26320 -6743 26392 -6728
use sky130_fd_pr__nfet_01v8_lvt_63HJ42  sky130_fd_pr__nfet_01v8_lvt_63HJ42_0
timestamp 1724943425
transform 1 0 19950 0 1 -9636
box -424 -257 424 257
use sky130_fd_pr__nfet_01v8_lvt_S7NVL3  sky130_fd_pr__nfet_01v8_lvt_S7NVL3_0
timestamp 1725190886
transform 1 0 19861 0 1 -8156
box -1883 -979 1883 979
use sky130_fd_pr__pfet_01v8_lvt_W4537V  sky130_fd_pr__pfet_01v8_lvt_W4537V_0
timestamp 1725004556
transform -1 0 22610 0 -1 -5723
box -1196 -973 1196 973
use sky130_fd_pr__pfet_01v8_lvt_WU9DQP  sky130_fd_pr__pfet_01v8_lvt_WU9DQP_0
timestamp 1725126992
transform 1 0 19872 0 1 -6222
box -323 -898 323 864
use sky130_fd_pr__res_xhigh_po_0p35_VRVSRL  sky130_fd_pr__res_xhigh_po_0p35_VRVSRL_0
timestamp 1724926688
transform -1 0 23753 0 -1 -8361
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p35_VUHUKX  sky130_fd_pr__res_xhigh_po_0p35_VUHUKX_0
timestamp 1725054279
transform -1 0 24547 0 -1 -8337
box -201 -672 201 672
use sky130_fd_pr__res_xhigh_po_0p35_Z5USRC  sky130_fd_pr__res_xhigh_po_0p35_Z5USRC_0
timestamp 1724926688
transform -1 0 25341 0 -1 -8361
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p69_5SXZXT  sky130_fd_pr__res_xhigh_po_0p69_5SXZXT_0
timestamp 1725054543
transform 1 0 24557 0 1 -9834
box -1522 -708 1522 708
use sky130_fd_pr__pfet_01v8_lvt_6GTY34  XM1
timestamp 1724939774
transform 1 0 25356 0 1 -5820
box -855 -1098 855 1064
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 5 1288
timestamp 1704896540
transform -1 0 33095 0 -1 -4445
box 0 0 1340 1340
<< labels >>
flabel metal1 26176 -8411 26288 -8297 0 FreeSans 160 0 0 0 Vbgr
port 2 nsew
flabel metal1 22344 -4599 22547 -4401 0 FreeSans 160 0 0 0 Vbgr
port 2 nsew
flabel metal3 20524 -4594 20654 -4534 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 22498 -7703 22598 -7591 0 FreeSans 160 0 0 0 VSS
port 3 nsew
flabel metal1 25949 -10812 26067 -10672 0 FreeSans 160 0 0 0 VSS
port 3 nsew
flabel metal1 19419 -9776 19489 -9658 0 FreeSans 160 0 0 0 VSS
port 3 nsew
rlabel metal1 19842 -9364 19900 -9306 1 Sop
rlabel metal2 20222 -7294 20326 -7200 1 PLUS
rlabel metal1 21102 -7155 21177 -7080 1 opout
rlabel metal2 23896 -7497 23996 -7397 1 MINUS
flabel space 23035 -12270 23165 -12097 0 FreeSans 160 0 0 0 VSS
port 3 nsew
rlabel metal1 20494 -9272 20576 -9210 1 Gcm2
rlabel metal1 20361 -9309 20495 -9175 1 Gcm2
flabel space 20395 -9810 20479 -9639 0 FreeSans 160 0 0 0 VSS
port 3 nsew
flabel space 22935 -6833 23044 -6780 0 FreeSans 160 0 0 0 VSS
port 3 nsew
flabel space 23031 -9138 23139 -9043 0 FreeSans 160 0 0 0 VSS
port 3 nsew
flabel metal1 16542 -7789 16772 -7510 0 FreeSans 160 0 0 0 VSS
port 3 nsew
rlabel metal2 19700 -5999 19799 -5798 1 Gcm1
<< end >>
