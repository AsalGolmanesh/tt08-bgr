** sch_path: /home/ttuser/tt08-bgr/xschem/core_PreL.sch
.subckt core_PreL MINUS PLUS Vbgr VDD VSS Vxy
*.PININFO MINUS:O PLUS:O Vbgr:O VDD:I VSS:I Vxy:I
XQ1 VSS VSS MINUS sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
XQ2 VSS VSS net1 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=33
XM1 MINUS Vxy VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XM2 PLUS Vxy VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XM3 Vbgr Vxy VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XR2 VSS net3 VSS sky130_fd_pr__res_xhigh_po W=1 L=11 mult=1 m=1
XR3 VSS net4 VSS sky130_fd_pr__res_xhigh_po W=1 L=11 mult=1 m=1
XR4 net2 Vbgr VSS sky130_fd_pr__res_xhigh_po W=1 L=12 mult=1 m=1
XR25 VSS net2 VSS sky130_fd_pr__res_xhigh_po W=1 L=12 mult=1 m=1
XR1 net1 net6 VSS sky130_fd_pr__res_xhigh_po W=1 L=1 mult=1 m=1
XR19 net3 PLUS VSS sky130_fd_pr__res_xhigh_po W=1 L=11 mult=1 m=1
XR21 net6 net5 VSS sky130_fd_pr__res_xhigh_po W=1 L=1 mult=1 m=1
XR22 net5 PLUS VSS sky130_fd_pr__res_xhigh_po W=1 L=1 mult=1 m=1
XR24 net4 MINUS net7 sky130_fd_pr__res_xhigh_po W=1 L=11 mult=1 m=1
.ends
.end
