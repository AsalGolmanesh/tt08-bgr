* NGSPICE file created from core_prel_parax.ext - technology: sky130A

.subckt core_prel_parax VDD Vbgr VSS
X0 VDD.t24 opout.t11 PLUS.t2 VDD.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 VSS.t76 VSS.t77 VSS.t75 sky130_fd_pr__res_xhigh_po_0p35 l=1
X2 a_24605_n9724# a_24371_n10376# VSS.t87 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X3 VSS.t78 Vbgr.t3 opout.t4 opout.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X4 Gcm2 opout.t12 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X5 MINUS.t3 opout.t13 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X6 VSS.t30 VSS.t27 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X7 VSS.t35 VSS.t64 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X8 VSS.t32 VSS.t63 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X9 VSS.t32 VSS.t62 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X10 a_23884_n8277# a_23718_n8877# VSS.t73 sky130_fd_pr__res_xhigh_po_0p35 l=1
X11 VSS.t35 VSS.t61 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X12 VSS.t32 VSS.t60 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X13 VSS.t32 VSS.t59 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X14 VDD.t18 opout.t14 Vbgr.t2 VDD.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X15 a_24137_n9724# a_23903_n10376# VSS.t74 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X16 VSS.t35 VSS.t58 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X17 VSS.t32 VSS.t57 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X18 VSS.t83 Vbgr.t4 opout.t8 opout.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X19 Sop MINUS.t4 opout.t0 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=4
X20 VSS.t32 VSS.t56 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X21 VDD.t1 Gcm1.t0 Gcm1.t1 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=1
X22 VSS.t17 VSS.t18 VSS.t16 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X23 VSS.t32 VSS.t55 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X24 VSS.t32 VSS.t65 MINUS.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X25 PLUS.t1 XQ2[0|0].Emitter VSS.t21 sky130_fd_pr__res_xhigh_po_0p35 l=0.9
X26 a_24974_n8277# a_24808_n8877# VSS.t66 sky130_fd_pr__res_xhigh_po_0p35 l=1
X27 a_24974_n8277# a_25472_n8877# VSS.t86 sky130_fd_pr__res_xhigh_po_0p35 l=1
X28 PLUS.t0 a_25472_n8877# VSS.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1
X29 VSS.t32 VSS.t54 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X30 VSS.t32 VSS.t53 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X31 Vbgr.t0 a_25307_n10376# VSS.t15 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X32 VSS.t81 VSS.t82 VSS.t80 sky130_fd_pr__res_xhigh_po_0p35 l=1
X33 a_23669_n9724# a_23435_n10376# VSS.t7 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X34 a_23669_n9724# a_23903_n10376# VSS.t85 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X35 VDD.t8 VDD.t6 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=0.5
X36 a_25073_n9724# a_24839_n10376# VSS.t26 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X37 VSS.t32 VSS.t52 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X38 VSS.t32 VSS.t51 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X39 VSS.t32 VSS.t50 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X40 VDD.t16 opout.t15 Gcm2 VDD.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X41 VDD.t14 opout.t16 MINUS.t2 VDD.t13 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X42 Sop PLUS.t4 Gcm1.t3 VSS.t71 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X43 Sop Gcm2 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X44 Gcm2 Gcm2 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X45 VSS.t32 VSS.t49 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X46 opout.t10 Gcm1.t4 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=1
X47 VSS.t24 a_23435_n10376# VSS.t23 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X48 VSS.t32 VSS.t48 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X49 VSS.t32 VSS.t47 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X50 VSS.t32 VSS.t46 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X51 VSS.t32 VSS.t45 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X52 VSS.t13 VSS.t14 VSS.t12 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X53 VSS.t35 VSS.t44 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X54 PLUS.t3 opout.t17 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X55 VSS.t32 VSS.t43 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X56 VDD.t5 VDD.t2 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.5
X57 a_25073_n9724# a_25307_n10376# VSS.t11 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X58 VSS.t90 a_23718_n8877# VSS.t89 sky130_fd_pr__res_xhigh_po_0p35 l=1
X59 VSS.t32 VSS.t42 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X60 VSS.t32 VSS.t41 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X61 a_23386_n8277# a_23552_n8877# VSS.t9 sky130_fd_pr__res_xhigh_po_0p35 l=1
X62 a_24050_n8277# a_24216_n8877# VSS.t10 sky130_fd_pr__res_xhigh_po_0p35 l=1
X63 a_24050_n8277# a_23552_n8877# VSS.t84 sky130_fd_pr__res_xhigh_po_0p35 l=1
X64 a_24137_n9724# a_24371_n10376# VSS.t6 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X65 Gcm1.t2 PLUS.t5 Sop VSS.t70 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=4
X66 VSS.t32 VSS.t40 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X67 Vbgr.t1 opout.t18 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X68 opout.t9 MINUS.t5 Sop VSS.t88 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X69 a_23884_n8277# a_24808_n8877# VSS.t72 sky130_fd_pr__res_xhigh_po_0p35 l=1
X70 VSS.t1 Gcm2 Sop VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X71 VSS.t39 VSS.t37 Gcm2 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X72 VSS.t32 VSS.t36 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X73 a_25140_n8277# a_24216_n8877# VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X74 a_25140_n8277# MINUS.t0 VSS.t22 sky130_fd_pr__res_xhigh_po_0p35 l=1
X75 a_24605_n9724# a_24839_n10376# VSS.t19 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X76 VSS.t35 VSS.t34 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X77 VSS.t67 Vbgr.t5 opout.t2 opout.t1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X78 VSS.t32 VSS.t33 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X79 VSS.t32 VSS.t31 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X80 VSS.t79 Vbgr.t6 opout.t6 opout.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X81 a_23386_n8277# VSS.t69 VSS.t68 sky130_fd_pr__res_xhigh_po_0p35 l=1
R0 opout.n1 opout.t14 674.212
R1 opout.n1 opout.t12 674.149
R2 opout.n1 opout.t15 674.149
R3 opout.n1 opout.t17 674.149
R4 opout.n1 opout.t11 674.149
R5 opout.n1 opout.t13 674.149
R6 opout.n1 opout.t16 674.149
R7 opout.n1 opout.t18 674.149
R8 opout.n4 opout.t10 232.543
R9 opout.n0 opout.t6 228.483
R10 opout.n0 opout.t2 228.215
R11 opout.n0 opout.t8 228.215
R12 opout.n0 opout.t4 228.215
R13 opout.n4 opout.n3 211.4
R14 opout.t1 opout.t5 173.161
R15 opout.t7 opout.t3 173.161
R16 opout.n2 opout.t1 86.5808
R17 opout.n2 opout.t7 86.5808
R18 opout.n0 opout.n2 16.5121
R19 opout.n0 opout.n1 8.29418
R20 opout.n3 opout.t0 2.1755
R21 opout.n3 opout.t9 2.1755
R22 opout.n4 opout.n0 1.94511
R23 PLUS.n2 PLUS.n0 276.264
R24 PLUS.n3 PLUS.t5 67.4131
R25 PLUS.n3 PLUS.t4 66.1779
R26 PLUS.n1 PLUS.t1 53.7169
R27 PLUS.n1 PLUS.t0 43.8915
R28 PLUS PLUS.n2 10.7127
R29 PLUS PLUS.n3 7.65631
R30 PLUS.n0 PLUS.t2 2.857
R31 PLUS.n0 PLUS.t3 2.857
R32 PLUS.n2 PLUS.n1 0.40761
R33 VDD.n2 VDD.t6 675.381
R34 VDD.n13 VDD.t2 674.89
R35 VDD.n21 VDD.t0 385.031
R36 VDD.n24 VDD.t25 374.053
R37 VDD.n15 VDD.t5 278.337
R38 VDD.t8 VDD.n1 278.334
R39 VDD.n12 VDD.n11 275.077
R40 VDD.n10 VDD.n9 275.077
R41 VDD.n8 VDD.n7 275.077
R42 VDD.n6 VDD.n5 275.077
R43 VDD.n4 VDD.n3 275.077
R44 VDD.n23 VDD.n22 227.799
R45 VDD.n18 VDD.n17 162.465
R46 VDD.n16 VDD.n14 152.345
R47 VDD.t3 VDD.n16 143.857
R48 VDD.n17 VDD.t7 140.78
R49 VDD.t0 VDD.t25 139.103
R50 VDD.n17 VDD.n1 118.692
R51 VDD.n16 VDD.n15 116.584
R52 VDD.t7 VDD.t17 69.427
R53 VDD.t17 VDD.t9 69.427
R54 VDD.t9 VDD.t13 69.427
R55 VDD.t13 VDD.t19 69.427
R56 VDD.t19 VDD.t23 69.427
R57 VDD.t23 VDD.t11 69.427
R58 VDD.t11 VDD.t15 69.427
R59 VDD.t15 VDD.t21 69.427
R60 VDD.t21 VDD.t3 69.427
R61 VDD.n22 VDD.t26 3.57113
R62 VDD.n22 VDD.t1 3.57113
R63 VDD.n11 VDD.t22 2.857
R64 VDD.n11 VDD.t4 2.857
R65 VDD.n9 VDD.t12 2.857
R66 VDD.n9 VDD.t16 2.857
R67 VDD.n7 VDD.t20 2.857
R68 VDD.n7 VDD.t24 2.857
R69 VDD.n5 VDD.t10 2.857
R70 VDD.n5 VDD.t14 2.857
R71 VDD.n3 VDD.t8 2.857
R72 VDD.n3 VDD.t18 2.857
R73 VDD.n14 VDD.n0 2.26217
R74 VDD.n19 VDD.n18 2.26217
R75 VDD.n19 VDD.n1 2.09911
R76 VDD.n15 VDD.n0 1.99684
R77 VDD.n21 VDD 1.32496
R78 VDD.n25 VDD.n24 1.29507
R79 VDD.n26 VDD.n20 0.975159
R80 VDD.n20 VDD.n19 0.723704
R81 VDD.n23 VDD.n21 0.286437
R82 VDD.n24 VDD.n23 0.275891
R83 VDD.n20 VDD.n0 0.218658
R84 VDD.n26 VDD.n25 0.214974
R85 VDD.n13 VDD.n12 0.143692
R86 VDD.n4 VDD.n2 0.1405
R87 VDD.n6 VDD.n4 0.122038
R88 VDD.n8 VDD.n6 0.122038
R89 VDD.n10 VDD.n8 0.122038
R90 VDD.n12 VDD.n10 0.122038
R91 VDD VDD.n26 0.04985
R92 VDD.n26 VDD 0.0299078
R93 VDD.n25 VDD 0.00829732
R94 VDD.n14 VDD.n13 0.00176918
R95 VDD.n18 VDD.n2 0.00165385
R96 VSS.n4313 VSS.n2055 122426
R97 VSS.n4304 VSS.n2055 35909.3
R98 VSS.n4311 VSS.n4232 15870.1
R99 VSS.n4291 VSS.n4238 12208.2
R100 VSS.n4278 VSS.n4277 7289
R101 VSS.n4279 VSS.n4277 7289
R102 VSS.n4263 VSS.n4254 7289
R103 VSS.n4264 VSS.n4254 7289
R104 VSS.n4255 VSS.n4249 6993.5
R105 VSS.n4269 VSS.n4250 6993.5
R106 VSS.n4318 VSS.n2055 6981.01
R107 VSS.n4335 VSS.n4318 4974.74
R108 VSS.n4279 VSS.n4269 3743
R109 VSS.n4264 VSS.n4255 3743
R110 VSS.n4278 VSS.n4250 3644.5
R111 VSS.n4263 VSS.n4249 3644.5
R112 VSS.n4335 VSS.n4334 3409.8
R113 VSS.t35 VSS.n1746 2890.74
R114 VSS.n4655 VSS.n1702 2277.04
R115 VSS.n4310 VSS.n4309 2062.31
R116 VSS.n3187 VSS.n3186 1851.56
R117 VSS.n4308 VSS.n4231 1679.57
R118 VSS.n2626 VSS.n2588 1634.59
R119 VSS.n2691 VSS.n2661 1559.06
R120 VSS.n2691 VSS.n2690 1559.06
R121 VSS.n2690 VSS.n2689 1559.06
R122 VSS.n2689 VSS.n2667 1559.06
R123 VSS.n2667 VSS.n1736 1559.06
R124 VSS.n2681 VSS.n1737 1559.06
R125 VSS.n2681 VSS.n2680 1559.06
R126 VSS.n2680 VSS.n2679 1559.06
R127 VSS.n2679 VSS.n2673 1559.06
R128 VSS.n2673 VSS.n1738 1559.06
R129 VSS.n3186 VSS.n3185 1559.06
R130 VSS.n3185 VSS.n3156 1559.06
R131 VSS.n3179 VSS.n3156 1559.06
R132 VSS.n3179 VSS.n3178 1559.06
R133 VSS.n3175 VSS.n3174 1559.06
R134 VSS.n3174 VSS.n3173 1559.06
R135 VSS.n3173 VSS.n3161 1559.06
R136 VSS.n3165 VSS.n3161 1559.06
R137 VSS.n3166 VSS.n3165 1559.06
R138 VSS.n4329 VSS.n4328 1540.86
R139 VSS.n4328 VSS.n4327 1540.86
R140 VSS.n4327 VSS.n1747 1540.86
R141 VSS.n4638 VSS.n1732 1540.86
R142 VSS.n4644 VSS.n1732 1540.86
R143 VSS.n4645 VSS.n4644 1540.86
R144 VSS.n4648 VSS.n4645 1540.86
R145 VSS.n4648 VSS.n4647 1540.86
R146 VSS.n4647 VSS.n4646 1540.86
R147 VSS.n4656 VSS.n4655 1540.86
R148 VSS.n4680 VSS.n4656 1540.86
R149 VSS.n4680 VSS.n4679 1540.86
R150 VSS.n4679 VSS.n4678 1540.86
R151 VSS.n4678 VSS.n4657 1540.86
R152 VSS.n4672 VSS.n4671 1540.86
R153 VSS.n4671 VSS.n4670 1540.86
R154 VSS.n4670 VSS.n4661 1540.86
R155 VSS.n4664 VSS.n4661 1540.86
R156 VSS.n4664 VSS.n4663 1540.86
R157 VSS.n4289 VSS.n4240 1332.39
R158 VSS.n4243 VSS.n4239 1311.29
R159 VSS.n4646 VSS.n1702 1284.05
R160 VSS.t35 VSS.n1736 1056.69
R161 VSS.n3178 VSS.t32 1056.69
R162 VSS.t35 VSS.n1747 1044.36
R163 VSS.n4657 VSS.t32 1044.36
R164 VSS.n4255 VSS.n4248 857.529
R165 VSS.n4269 VSS.n4248 857.529
R166 VSS.n2598 VSS.n1702 855.557
R167 VSS.n4038 VSS.t32 855.557
R168 VSS.n4065 VSS.t32 855.557
R169 VSS.n4081 VSS.n4075 855.557
R170 VSS.n4099 VSS.n4091 855.557
R171 VSS.n4284 VSS.n4249 840.148
R172 VSS.n4284 VSS.n4250 840.148
R173 VSS.n4317 VSS.n4229 827.635
R174 VSS.n4317 VSS.n4316 785.924
R175 VSS.n4247 VSS.n4229 766.952
R176 VSS.n4336 VSS.n4335 728.679
R177 VSS.n4287 VSS.n4230 724.09
R178 VSS.n4334 VSS.n4319 718.693
R179 VSS.n3098 VSS.n3097 665.731
R180 VSS.t35 VSS.n1740 665.731
R181 VSS.t35 VSS.n1753 665.731
R182 VSS.t35 VSS.n1750 665.731
R183 VSS.t35 VSS.n1738 658.269
R184 VSS.n3166 VSS.t32 658.269
R185 VSS.n3097 VSS.n3096 648.096
R186 VSS.t35 VSS.n1739 648.096
R187 VSS.t35 VSS.n4637 648.096
R188 VSS.t35 VSS.n1751 648.096
R189 VSS.n4191 VSS.n4156 641.164
R190 VSS.n4663 VSS.n1245 616.342
R191 VSS.n5350 VSS.n194 585
R192 VSS.n5350 VSS.n5349 585
R193 VSS.n218 VSS.n202 585
R194 VSS.n5344 VSS.n218 585
R195 VSS.n3634 VSS.n220 585
R196 VSS.n5006 VSS.n5005 585
R197 VSS.n5026 VSS.n699 585
R198 VSS.n5027 VSS.n5026 585
R199 VSS.n4841 VSS.n186 585
R200 VSS.n5360 VSS.n186 585
R201 VSS.n4841 VSS.n187 585
R202 VSS.n5360 VSS.n187 585
R203 VSS.n5032 VSS.n185 585
R204 VSS.n5360 VSS.n185 585
R205 VSS.n5032 VSS.n188 585
R206 VSS.n5360 VSS.n188 585
R207 VSS.n5358 VSS.n184 585
R208 VSS.n5360 VSS.n184 585
R209 VSS.n5359 VSS.n5358 585
R210 VSS.n5360 VSS.n5359 585
R211 VSS.n4197 VSS.n69 585
R212 VSS.n5357 VSS.n189 585
R213 VSS.n5357 VSS.n5356 585
R214 VSS.n5031 VSS.n693 585
R215 VSS.n5031 VSS.n5030 585
R216 VSS.n4840 VSS.n886 585
R217 VSS.n4840 VSS.n4839 585
R218 VSS.n4839 VSS.n69 585
R219 VSS.n4839 VSS.n888 585
R220 VSS.n888 VSS.n886 585
R221 VSS.n886 VSS.n71 585
R222 VSS.n5030 VSS.n5029 585
R223 VSS.n5030 VSS.n71 585
R224 VSS.n5029 VSS.n693 585
R225 VSS.n693 VSS.n71 585
R226 VSS.n5356 VSS.n5355 585
R227 VSS.n5356 VSS.n71 585
R228 VSS.n5355 VSS.n189 585
R229 VSS.n189 VSS.n71 585
R230 VSS.n996 VSS.n995 585
R231 VSS.n995 VSS.n994 585
R232 VSS.n1033 VSS.n998 585
R233 VSS.n958 VSS.n225 585
R234 VSS.n5341 VSS.n225 585
R235 VSS.n958 VSS.n226 585
R236 VSS.n5341 VSS.n226 585
R237 VSS.n5011 VSS.n224 585
R238 VSS.n5341 VSS.n224 585
R239 VSS.n5011 VSS.n227 585
R240 VSS.n5341 VSS.n227 585
R241 VSS.n5342 VSS.n219 585
R242 VSS.n5342 VSS.n5341 585
R243 VSS.n221 VSS.n219 585
R244 VSS.n5341 VSS.n221 585
R245 VSS.n4097 VSS.n27 585
R246 VSS.n3805 VSS.n3631 585
R247 VSS.n3631 VSS.n222 585
R248 VSS.n5010 VSS.n718 585
R249 VSS.n5010 VSS.n5009 585
R250 VSS.n1177 VSS.n955 585
R251 VSS.n1179 VSS.n955 585
R252 VSS.n1179 VSS.n27 585
R253 VSS.n1179 VSS.n1178 585
R254 VSS.n1178 VSS.n1177 585
R255 VSS.n1177 VSS.n29 585
R256 VSS.n5009 VSS.n5008 585
R257 VSS.n5009 VSS.n29 585
R258 VSS.n5008 VSS.n718 585
R259 VSS.n718 VSS.n29 585
R260 VSS.n3806 VSS.n222 585
R261 VSS.n222 VSS.n29 585
R262 VSS.n3806 VSS.n3805 585
R263 VSS.n3805 VSS.n29 585
R264 VSS.n607 VSS.n575 585
R265 VSS.n5339 VSS.n223 585
R266 VSS.n5341 VSS.n223 585
R267 VSS.n5340 VSS.n5339 585
R268 VSS.n5341 VSS.n5340 585
R269 VSS.n5338 VSS.n228 585
R270 VSS.n228 VSS.n27 585
R271 VSS.n5338 VSS.n5337 585
R272 VSS.n5337 VSS.n5336 585
R273 VSS.n5337 VSS.n29 585
R274 VSS.n5336 VSS.n228 585
R275 VSS.n5334 VSS.n5333 585
R276 VSS.n5362 VSS.n180 585
R277 VSS.n5360 VSS.n180 585
R278 VSS.n5362 VSS.n5361 585
R279 VSS.n5361 VSS.n5360 585
R280 VSS.n182 VSS.n181 585
R281 VSS.n182 VSS.n69 585
R282 VSS.n572 VSS.n181 585
R283 VSS.n610 VSS.n572 585
R284 VSS.n572 VSS.n71 585
R285 VSS.n610 VSS.n182 585
R286 VSS.n608 VSS.n607 585
R287 VSS.n5377 VSS.n163 585
R288 VSS.n5047 VSS.n676 585
R289 VSS.n4856 VSS.n869 585
R290 VSS.n2206 VSS.n2205 585
R291 VSS.n3418 VSS.n3417 585
R292 VSS.n3954 VSS.n3922 585
R293 VSS.n5084 VSS.n5054 585
R294 VSS.n4560 VSS.n4559 585
R295 VSS.n2998 VSS.n2965 585
R296 VSS.n2963 VSS.n2930 585
R297 VSS.n1954 VSS.n1952 585
R298 VSS.n3961 VSS.n1952 585
R299 VSS.n1954 VSS.n1890 585
R300 VSS.n3961 VSS.n1890 585
R301 VSS.n2983 VSS.n2211 585
R302 VSS.n3961 VSS.n2211 585
R303 VSS.n2983 VSS.n2213 585
R304 VSS.n3961 VSS.n2213 585
R305 VSS.n3959 VSS.n2210 585
R306 VSS.n3961 VSS.n2210 585
R307 VSS.n3960 VSS.n3959 585
R308 VSS.n3961 VSS.n3960 585
R309 VSS.n2209 VSS.n2208 585
R310 VSS.n3961 VSS.n2209 585
R311 VSS.n3962 VSS.n2208 585
R312 VSS.n3962 VSS.n3961 585
R313 VSS.n2114 VSS.n2067 585
R314 VSS.n3963 VSS.n2170 585
R315 VSS.n2171 VSS.n2170 585
R316 VSS.n3958 VSS.n2214 585
R317 VSS.n3958 VSS.n3957 585
R318 VSS.n3443 VSS.n2325 585
R319 VSS.n2329 VSS.n2325 585
R320 VSS.n4563 VSS.n1889 585
R321 VSS.n1950 VSS.n1889 585
R322 VSS.n4780 VSS.n1250 585
R323 VSS.n1252 VSS.n1250 585
R324 VSS.n1844 VSS.n1250 585
R325 VSS.n4562 VSS.n1950 585
R326 VSS.n1950 VSS.n1844 585
R327 VSS.n4563 VSS.n4562 585
R328 VSS.n4563 VSS.n1844 585
R329 VSS.n3444 VSS.n2329 585
R330 VSS.n2329 VSS.n1844 585
R331 VSS.n3444 VSS.n3443 585
R332 VSS.n3443 VSS.n1844 585
R333 VSS.n3957 VSS.n3956 585
R334 VSS.n3957 VSS.n1844 585
R335 VSS.n3956 VSS.n2214 585
R336 VSS.n2214 VSS.n1844 585
R337 VSS.n3964 VSS.n2171 585
R338 VSS.n2171 VSS.n1844 585
R339 VSS.n3964 VSS.n3963 585
R340 VSS.n3963 VSS.n1844 585
R341 VSS.n2067 VSS.n2065 585
R342 VSS.n2067 VSS.n1844 585
R343 VSS.n4526 VSS.n4525 585
R344 VSS.n2697 VSS.n2692 585
R345 VSS.n2697 VSS.n2696 585
R346 VSS.n3061 VSS.n2748 585
R347 VSS.n3059 VSS.n2748 585
R348 VSS.n3061 VSS.n3060 585
R349 VSS.n3060 VSS.n3059 585
R350 VSS.n3060 VSS.n1748 585
R351 VSS.n3026 VSS.n2810 585
R352 VSS.n2810 VSS.n1757 585
R353 VSS.n3026 VSS.n3025 585
R354 VSS.n3025 VSS.n1757 585
R355 VSS.n3025 VSS.n1744 585
R356 VSS.n4498 VSS.n1998 585
R357 VSS.n4498 VSS.n4497 585
R358 VSS.n4496 VSS.n1998 585
R359 VSS.n4497 VSS.n4496 585
R360 VSS.n4496 VSS.n1745 585
R361 VSS.n3154 VSS.n2496 585
R362 VSS.n3188 VSS.n2496 585
R363 VSS.n3386 VSS.n2461 585
R364 VSS.n3420 VSS.n2461 585
R365 VSS.n2461 VSS.n1748 585
R366 VSS.n3001 VSS.n2903 585
R367 VSS.n3001 VSS.n3000 585
R368 VSS.n3001 VSS.n1744 585
R369 VSS.n4521 VSS.n1965 585
R370 VSS.n4523 VSS.n4521 585
R371 VSS.n4521 VSS.n1745 585
R372 VSS.n4523 VSS.n4522 585
R373 VSS.n4522 VSS.n1672 585
R374 VSS.n1965 VSS.n1964 585
R375 VSS.n1964 VSS.n1672 585
R376 VSS.n3000 VSS.n2928 585
R377 VSS.n2928 VSS.n1672 585
R378 VSS.n2904 VSS.n2903 585
R379 VSS.n2904 VSS.n1672 585
R380 VSS.n3420 VSS.n2462 585
R381 VSS.n2462 VSS.n1672 585
R382 VSS.n3386 VSS.n3385 585
R383 VSS.n3385 VSS.n1672 585
R384 VSS.n3188 VSS.n2497 585
R385 VSS.n2497 VSS.n1672 585
R386 VSS.n3154 VSS.n3153 585
R387 VSS.n3153 VSS.n1672 585
R388 VSS.n4687 VSS.n1701 585
R389 VSS.n4687 VSS.n1703 585
R390 VSS.n4687 VSS.n1695 585
R391 VSS.n4687 VSS.n1704 585
R392 VSS.n4687 VSS.n1689 585
R393 VSS.n4687 VSS.n1705 585
R394 VSS.n4687 VSS.n1683 585
R395 VSS.n4687 VSS.n1706 585
R396 VSS.n4687 VSS.n1677 585
R397 VSS.n4687 VSS.n4686 585
R398 VSS.n3188 VSS.n2495 585
R399 VSS.n3188 VSS.n3187 585
R400 VSS.n3386 VSS.n2460 585
R401 VSS.n3420 VSS.n2460 585
R402 VSS.n3419 VSS.n3386 585
R403 VSS.n3420 VSS.n3419 585
R404 VSS.n3419 VSS.n3418 585
R405 VSS.n2907 VSS.n2903 585
R406 VSS.n3000 VSS.n2907 585
R407 VSS.n2999 VSS.n2903 585
R408 VSS.n3000 VSS.n2999 585
R409 VSS.n2999 VSS.n2998 585
R410 VSS.n1990 VSS.n1965 585
R411 VSS.n4523 VSS.n1990 585
R412 VSS.n4524 VSS.n1965 585
R413 VSS.n4524 VSS.n4523 585
R414 VSS.n4525 VSS.n4524 585
R415 VSS.n5379 VSS.n158 585
R416 VSS.n162 VSS.n158 585
R417 VSS.n2205 VSS.n158 585
R418 VSS.n5086 VSS.n658 585
R419 VSS.n3922 VSS.n658 585
R420 VSS.n5053 VSS.n658 585
R421 VSS.n5049 VSS.n672 585
R422 VSS.n2930 VSS.n672 585
R423 VSS.n675 VSS.n672 585
R424 VSS.n4858 VSS.n864 585
R425 VSS.n868 VSS.n864 585
R426 VSS.n4559 VSS.n864 585
R427 VSS.n868 VSS.n665 585
R428 VSS.n5051 VSS.n665 585
R429 VSS.n4858 VSS.n667 585
R430 VSS.n5051 VSS.n667 585
R431 VSS.n675 VSS.n664 585
R432 VSS.n5051 VSS.n664 585
R433 VSS.n5050 VSS.n5049 585
R434 VSS.n5051 VSS.n5050 585
R435 VSS.n5053 VSS.n5052 585
R436 VSS.n5052 VSS.n5051 585
R437 VSS.n5086 VSS.n656 585
R438 VSS.n5051 VSS.n656 585
R439 VSS.n630 VSS.n162 585
R440 VSS.n5051 VSS.n630 585
R441 VSS.n5379 VSS.n156 585
R442 VSS.n5051 VSS.n156 585
R443 VSS.n5413 VSS.n129 585
R444 VSS.n5381 VSS.n129 585
R445 VSS.n5120 VSS.n129 585
R446 VSS.n5088 VSS.n129 585
R447 VSS.n663 VSS.n129 585
R448 VSS.n668 VSS.n129 585
R449 VSS.n4892 VSS.n129 585
R450 VSS.n4860 VSS.n129 585
R451 VSS.n4739 VSS.n129 585
R452 VSS.n1484 VSS.n129 585
R453 VSS.n5379 VSS.n157 585
R454 VSS.n162 VSS.n157 585
R455 VSS.n5379 VSS.n5378 585
R456 VSS.n5378 VSS.n162 585
R457 VSS.n5378 VSS.n5377 585
R458 VSS.n5086 VSS.n657 585
R459 VSS.n5053 VSS.n657 585
R460 VSS.n5086 VSS.n5085 585
R461 VSS.n5085 VSS.n5053 585
R462 VSS.n5085 VSS.n5084 585
R463 VSS.n5049 VSS.n671 585
R464 VSS.n675 VSS.n671 585
R465 VSS.n5049 VSS.n5048 585
R466 VSS.n5048 VSS.n675 585
R467 VSS.n5048 VSS.n5047 585
R468 VSS.n4858 VSS.n863 585
R469 VSS.n868 VSS.n863 585
R470 VSS.n4858 VSS.n4857 585
R471 VSS.n4857 VSS.n868 585
R472 VSS.n4857 VSS.n4856 585
R473 VSS.n1509 VSS.n1386 585
R474 VSS.n1386 VSS.n69 585
R475 VSS.n1386 VSS.n1383 585
R476 VSS.n1557 VSS.n1381 585
R477 VSS.n1557 VSS.n27 585
R478 VSS.n1557 VSS.n1556 585
R479 VSS.n5332 VSS.n5331 585
R480 VSS.n5333 VSS.n5332 585
R481 VSS.n3646 VSS.n3634 585
R482 VSS.n3646 VSS.n312 585
R483 VSS.n5004 VSS.n293 585
R484 VSS.n5005 VSS.n5004 585
R485 VSS.n1006 VSS.n998 585
R486 VSS.n1006 VSS.n273 585
R487 VSS.n5328 VSS.n273 585
R488 VSS.n293 VSS.n271 585
R489 VSS.n312 VSS.n270 585
R490 VSS.n5331 VSS.n5330 585
R491 VSS.n5329 VSS.n12 585
R492 VSS.n5499 VSS.n5498 585
R493 VSS.n5501 VSS.n11 585
R494 VSS.n5504 VSS.n5503 585
R495 VSS.n8 VSS.n7 585
R496 VSS.n5511 VSS.n5510 585
R497 VSS.n5514 VSS.n5513 585
R498 VSS.n5 VSS.n0 585
R499 VSS.n485 VSS.n1 585
R500 VSS.n489 VSS.n488 585
R501 VSS.n491 VSS.n482 585
R502 VSS.n497 VSS.n496 585
R503 VSS.n494 VSS.n493 585
R504 VSS.n327 VSS.n268 585
R505 VSS.n330 VSS.n329 585
R506 VSS.n5201 VSS.n5200 585
R507 VSS.n5203 VSS.n326 585
R508 VSS.n5206 VSS.n5205 585
R509 VSS.n323 VSS.n322 585
R510 VSS.n5216 VSS.n5215 585
R511 VSS.n5218 VSS.n321 585
R512 VSS.n5221 VSS.n5220 585
R513 VSS.n318 VSS.n314 585
R514 VSS.n5232 VSS.n5231 585
R515 VSS.n5234 VSS.n313 585
R516 VSS.n5238 VSS.n5237 585
R517 VSS.n309 VSS.n308 585
R518 VSS.n5247 VSS.n5246 585
R519 VSS.n5249 VSS.n307 585
R520 VSS.n5252 VSS.n5251 585
R521 VSS.n304 VSS.n303 585
R522 VSS.n5262 VSS.n5261 585
R523 VSS.n5264 VSS.n302 585
R524 VSS.n5267 VSS.n5266 585
R525 VSS.n299 VSS.n295 585
R526 VSS.n5278 VSS.n5277 585
R527 VSS.n5280 VSS.n294 585
R528 VSS.n5284 VSS.n5283 585
R529 VSS.n290 VSS.n289 585
R530 VSS.n5293 VSS.n5292 585
R531 VSS.n5295 VSS.n288 585
R532 VSS.n5298 VSS.n5297 585
R533 VSS.n285 VSS.n284 585
R534 VSS.n5308 VSS.n5307 585
R535 VSS.n5310 VSS.n283 585
R536 VSS.n5313 VSS.n5312 585
R537 VSS.n280 VSS.n276 585
R538 VSS.n5324 VSS.n5323 585
R539 VSS.n5326 VSS.n275 585
R540 VSS.n1202 VSS.n274 585
R541 VSS.n1207 VSS.n1204 585
R542 VSS.n4818 VSS.n4817 585
R543 VSS.n4815 VSS.n4814 585
R544 VSS.n4811 VSS.n1208 585
R545 VSS.n1211 VSS.n1209 585
R546 VSS.n4806 VSS.n4805 585
R547 VSS.n4803 VSS.n4802 585
R548 VSS.n4798 VSS.n1212 585
R549 VSS.n1217 VSS.n1214 585
R550 VSS.n4793 VSS.n4792 585
R551 VSS.n4790 VSS.n4789 585
R552 VSS.n2589 VSS.n2588 585
R553 VSS.n2621 VSS.n2620 585
R554 VSS.n2591 VSS.n2590 585
R555 VSS.n2619 VSS.n2591 585
R556 VSS.n2617 VSS.n2616 585
R557 VSS.n2618 VSS.n2617 585
R558 VSS.n2615 VSS.n2593 585
R559 VSS.n2593 VSS.n2592 585
R560 VSS.n2614 VSS.n2613 585
R561 VSS.n2613 VSS.n1742 585
R562 VSS.n2612 VSS.n2594 585
R563 VSS.n2612 VSS.n1741 585
R564 VSS.n2611 VSS.n2596 585
R565 VSS.n2611 VSS.n2610 585
R566 VSS.n2605 VSS.n2595 585
R567 VSS.n2609 VSS.n2595 585
R568 VSS.n2607 VSS.n2606 585
R569 VSS.n2608 VSS.n2607 585
R570 VSS.n2604 VSS.n2078 585
R571 VSS.n2604 VSS.n2597 585
R572 VSS.n2603 VSS.n2602 585
R573 VSS.n2601 VSS.n2600 585
R574 VSS.n2599 VSS.n2598 585
R575 VSS.n2077 VSS.n2076 585
R576 VSS.n4015 VSS.n4014 585
R577 VSS.n4016 VSS.n4015 585
R578 VSS.n2075 VSS.n2074 585
R579 VSS.n4017 VSS.n2075 585
R580 VSS.n4021 VSS.n4020 585
R581 VSS.n4020 VSS.n4019 585
R582 VSS.n4022 VSS.n2073 585
R583 VSS.n4018 VSS.n2073 585
R584 VSS.n4024 VSS.n4023 585
R585 VSS.n4025 VSS.n4024 585
R586 VSS.n2072 VSS.n2071 585
R587 VSS.n4026 VSS.n2072 585
R588 VSS.n4029 VSS.n4028 585
R589 VSS.n4028 VSS.n4027 585
R590 VSS.n4030 VSS.n2070 585
R591 VSS.n2070 VSS.n2069 585
R592 VSS.n4033 VSS.n4032 585
R593 VSS.n4034 VSS.n4033 585
R594 VSS.n4031 VSS.n2066 585
R595 VSS.n4035 VSS.n2066 585
R596 VSS.n4037 VSS.n2068 585
R597 VSS.n4037 VSS.n4036 585
R598 VSS.n4040 VSS.n4039 585
R599 VSS.n4039 VSS.n4038 585
R600 VSS.n4041 VSS.n2064 585
R601 VSS.n2064 VSS.n2063 585
R602 VSS.n4043 VSS.n4042 585
R603 VSS.n4044 VSS.n4043 585
R604 VSS.n2062 VSS.n2061 585
R605 VSS.n4045 VSS.n2062 585
R606 VSS.n4049 VSS.n4048 585
R607 VSS.n4048 VSS.n4047 585
R608 VSS.n4050 VSS.n2060 585
R609 VSS.n4046 VSS.n2060 585
R610 VSS.n4052 VSS.n4051 585
R611 VSS.n4053 VSS.n4052 585
R612 VSS.n2059 VSS.n2058 585
R613 VSS.n4054 VSS.n2059 585
R614 VSS.n4058 VSS.n4057 585
R615 VSS.n4057 VSS.n4056 585
R616 VSS.n4059 VSS.n2057 585
R617 VSS.n4055 VSS.n2057 585
R618 VSS.n4223 VSS.n4222 585
R619 VSS.n4223 VSS.n2056 585
R620 VSS.n4226 VSS.n4225 585
R621 VSS.n4227 VSS.n128 585
R622 VSS.n4065 VSS.n4064 585
R623 VSS.n4066 VSS.n4061 585
R624 VSS.n4220 VSS.n4219 585
R625 VSS.n4219 VSS.n4218 585
R626 VSS.n4062 VSS.n4060 585
R627 VSS.n4217 VSS.n4062 585
R628 VSS.n4215 VSS.n4214 585
R629 VSS.n4216 VSS.n4215 585
R630 VSS.n4213 VSS.n4068 585
R631 VSS.n4068 VSS.n4067 585
R632 VSS.n4212 VSS.n4211 585
R633 VSS.n4211 VSS.n4210 585
R634 VSS.n4070 VSS.n4069 585
R635 VSS.n4209 VSS.n4070 585
R636 VSS.n4207 VSS.n4206 585
R637 VSS.n4208 VSS.n4207 585
R638 VSS.n4205 VSS.n4072 585
R639 VSS.n4072 VSS.n4071 585
R640 VSS.n4204 VSS.n4203 585
R641 VSS.n4203 VSS.n4202 585
R642 VSS.n4201 VSS.n4074 585
R643 VSS.n4200 VSS.n4199 585
R644 VSS.n4081 VSS.n4076 585
R645 VSS.n4082 VSS.n4079 585
R646 VSS.n4156 VSS.n4155 585
R647 VSS.n4155 VSS.n4154 585
R648 VSS.n4080 VSS.n4077 585
R649 VSS.n4153 VSS.n4080 585
R650 VSS.n4151 VSS.n4150 585
R651 VSS.n4152 VSS.n4151 585
R652 VSS.n4149 VSS.n4084 585
R653 VSS.n4084 VSS.n4083 585
R654 VSS.n4148 VSS.n4147 585
R655 VSS.n4147 VSS.n4146 585
R656 VSS.n4086 VSS.n4085 585
R657 VSS.n4145 VSS.n4086 585
R658 VSS.n4143 VSS.n4142 585
R659 VSS.n4144 VSS.n4143 585
R660 VSS.n4141 VSS.n4088 585
R661 VSS.n4088 VSS.n4087 585
R662 VSS.n4140 VSS.n4139 585
R663 VSS.n4139 VSS.n4138 585
R664 VSS.n4137 VSS.n4090 585
R665 VSS.n4136 VSS.n4135 585
R666 VSS.n4099 VSS.n4092 585
R667 VSS.n4130 VSS.n4129 585
R668 VSS.n4102 VSS.n4098 585
R669 VSS.n4128 VSS.n4098 585
R670 VSS.n4126 VSS.n4125 585
R671 VSS.n4127 VSS.n4126 585
R672 VSS.n4124 VSS.n4101 585
R673 VSS.n4101 VSS.n4100 585
R674 VSS.n4123 VSS.n4122 585
R675 VSS.n4122 VSS.n4121 585
R676 VSS.n4120 VSS.n4103 585
R677 VSS.n4120 VSS.n4119 585
R678 VSS.n4107 VSS.n4104 585
R679 VSS.n4118 VSS.n4104 585
R680 VSS.n4116 VSS.n4115 585
R681 VSS.n4117 VSS.n4116 585
R682 VSS.n4114 VSS.n4106 585
R683 VSS.n4106 VSS.n4105 585
R684 VSS.n4113 VSS.n4112 585
R685 VSS.n4112 VSS.n4111 585
R686 VSS.n4110 VSS.n4109 585
R687 VSS.n4320 VSS.n2054 585
R688 VSS.n4336 VSS.n2054 585
R689 VSS.n4339 VSS.n4338 585
R690 VSS.n4338 VSS.n4337 585
R691 VSS.n4341 VSS.n2030 585
R692 VSS.n2030 VSS.n2029 585
R693 VSS.n4345 VSS.n4344 585
R694 VSS.n4346 VSS.n4345 585
R695 VSS.n2031 VSS.n2027 585
R696 VSS.n4347 VSS.n2027 585
R697 VSS.n4350 VSS.n4349 585
R698 VSS.n4349 VSS.n4348 585
R699 VSS.n2026 VSS.n2024 585
R700 VSS.n2028 VSS.n2026 585
R701 VSS.n4355 VSS.n2004 585
R702 VSS.n2004 VSS.n2003 585
R703 VSS.n4360 VSS.n4359 585
R704 VSS.n4361 VSS.n4360 585
R705 VSS.n2022 VSS.n2001 585
R706 VSS.n4362 VSS.n2001 585
R707 VSS.n4364 VSS.n2002 585
R708 VSS.n4364 VSS.n4363 585
R709 VSS.n4365 VSS.n2000 585
R710 VSS.n4365 VSS.n1751 585
R711 VSS.n4494 VSS.n4493 585
R712 VSS.n4494 VSS.n1750 585
R713 VSS.n4491 VSS.n4366 585
R714 VSS.n4486 VSS.n4366 585
R715 VSS.n4489 VSS.n4488 585
R716 VSS.n4488 VSS.n4487 585
R717 VSS.n4478 VSS.n4455 585
R718 VSS.n4485 VSS.n4455 585
R719 VSS.n4483 VSS.n4482 585
R720 VSS.n4484 VSS.n4483 585
R721 VSS.n4476 VSS.n4457 585
R722 VSS.n4457 VSS.n4456 585
R723 VSS.n4464 VSS.n4458 585
R724 VSS.n4468 VSS.n4464 585
R725 VSS.n4471 VSS.n4470 585
R726 VSS.n4470 VSS.n4469 585
R727 VSS.n4463 VSS.n4462 585
R728 VSS.n4467 VSS.n4463 585
R729 VSS.n4465 VSS.n1759 585
R730 VSS.n4466 VSS.n4465 585
R731 VSS.n4633 VSS.n1756 585
R732 VSS.n1756 VSS.n1754 585
R733 VSS.n4636 VSS.n4635 585
R734 VSS.n4637 VSS.n4636 585
R735 VSS.n3028 VSS.n3027 585
R736 VSS.n3028 VSS.n1753 585
R737 VSS.n3031 VSS.n3030 585
R738 VSS.n3030 VSS.n3029 585
R739 VSS.n3033 VSS.n2804 585
R740 VSS.n2804 VSS.n2803 585
R741 VSS.n3037 VSS.n3036 585
R742 VSS.n3038 VSS.n3037 585
R743 VSS.n2805 VSS.n2801 585
R744 VSS.n3039 VSS.n2801 585
R745 VSS.n3042 VSS.n3041 585
R746 VSS.n3041 VSS.n3040 585
R747 VSS.n2800 VSS.n2798 585
R748 VSS.n2802 VSS.n2800 585
R749 VSS.n3047 VSS.n2783 585
R750 VSS.n2783 VSS.n2782 585
R751 VSS.n3052 VSS.n3051 585
R752 VSS.n3053 VSS.n3052 585
R753 VSS.n2796 VSS.n2780 585
R754 VSS.n3054 VSS.n2780 585
R755 VSS.n3056 VSS.n2781 585
R756 VSS.n3056 VSS.n3055 585
R757 VSS.n3058 VSS.n3057 585
R758 VSS.n3057 VSS.n1739 585
R759 VSS.n3063 VSS.n3062 585
R760 VSS.n3063 VSS.n1740 585
R761 VSS.n3066 VSS.n3065 585
R762 VSS.n3065 VSS.n3064 585
R763 VSS.n3068 VSS.n2725 585
R764 VSS.n2725 VSS.n2724 585
R765 VSS.n3072 VSS.n3071 585
R766 VSS.n3073 VSS.n3072 585
R767 VSS.n2726 VSS.n2723 585
R768 VSS.n3074 VSS.n2723 585
R769 VSS.n3077 VSS.n3076 585
R770 VSS.n3076 VSS.n3075 585
R771 VSS.n2721 VSS.n2716 585
R772 VSS.n2716 VSS.n2715 585
R773 VSS.n3083 VSS.n3082 585
R774 VSS.n3084 VSS.n3083 585
R775 VSS.n2717 VSS.n2714 585
R776 VSS.n3085 VSS.n2714 585
R777 VSS.n3088 VSS.n3087 585
R778 VSS.n3087 VSS.n3086 585
R779 VSS.n3092 VSS.n2664 585
R780 VSS.n2664 VSS.n2662 585
R781 VSS.n3095 VSS.n3094 585
R782 VSS.n3096 VSS.n3095 585
R783 VSS.n2693 VSS.n2660 585
R784 VSS.n3098 VSS.n2660 585
R785 VSS.n3101 VSS.n3100 585
R786 VSS.n3100 VSS.n3099 585
R787 VSS.n3103 VSS.n2638 585
R788 VSS.n2638 VSS.n2637 585
R789 VSS.n3107 VSS.n3106 585
R790 VSS.n3108 VSS.n3107 585
R791 VSS.n2639 VSS.n2636 585
R792 VSS.n3109 VSS.n2636 585
R793 VSS.n3112 VSS.n3111 585
R794 VSS.n3111 VSS.n3110 585
R795 VSS.n2634 VSS.n2629 585
R796 VSS.n2629 VSS.n2628 585
R797 VSS.n3118 VSS.n3117 585
R798 VSS.n3119 VSS.n3118 585
R799 VSS.n2630 VSS.n2587 585
R800 VSS.n3120 VSS.n2587 585
R801 VSS.n3123 VSS.n3122 585
R802 VSS.n3122 VSS.n3121 585
R803 VSS.n2586 VSS.n2584 585
R804 VSS.n2627 VSS.n2586 585
R805 VSS.n2625 VSS.n2624 585
R806 VSS.n2626 VSS.n2625 585
R807 VSS.n4331 VSS.n4319 585
R808 VSS.n4334 VSS.n4333 585
R809 VSS.n4647 VSS.n1731 585
R810 VSS.n4650 VSS.n4649 585
R811 VSS.n4649 VSS.n4648 585
R812 VSS.n1730 VSS.n1729 585
R813 VSS.n4645 VSS.n1730 585
R814 VSS.n4643 VSS.n4642 585
R815 VSS.n4644 VSS.n4643 585
R816 VSS.n4641 VSS.n1733 585
R817 VSS.n1733 VSS.n1732 585
R818 VSS.n4640 VSS.n4639 585
R819 VSS.n4639 VSS.n4638 585
R820 VSS.n1735 VSS.n1734 585
R821 VSS.n1747 VSS.n1735 585
R822 VSS.n4326 VSS.n4325 585
R823 VSS.n4327 VSS.n4326 585
R824 VSS.n4324 VSS.n4322 585
R825 VSS.n4328 VSS.n4322 585
R826 VSS.n4330 VSS.n4323 585
R827 VSS.n4330 VSS.n4329 585
R828 VSS.n4646 VSS.n1708 585
R829 VSS.n1251 VSS.n1249 585
R830 VSS.n4663 VSS.n1249 585
R831 VSS.n4666 VSS.n4665 585
R832 VSS.n4665 VSS.n4664 585
R833 VSS.n4667 VSS.n4662 585
R834 VSS.n4662 VSS.n4661 585
R835 VSS.n4669 VSS.n4668 585
R836 VSS.n4670 VSS.n4669 585
R837 VSS.n4660 VSS.n4659 585
R838 VSS.n4671 VSS.n4660 585
R839 VSS.n4674 VSS.n4673 585
R840 VSS.n4673 VSS.n4672 585
R841 VSS.n4675 VSS.n4658 585
R842 VSS.n4658 VSS.n4657 585
R843 VSS.n4677 VSS.n4676 585
R844 VSS.n4678 VSS.n4677 585
R845 VSS.n4653 VSS.n4651 585
R846 VSS.n4679 VSS.n4653 585
R847 VSS.n4682 VSS.n4681 585
R848 VSS.n4681 VSS.n4680 585
R849 VSS.n4656 VSS.n4652 585
R850 VSS.n4655 VSS.n4654 585
R851 VSS.n4782 VSS.n4781 585
R852 VSS.n1406 VSS.n1405 585
R853 VSS.n1404 VSS.n1403 585
R854 VSS.n1402 VSS.n1401 585
R855 VSS.n1400 VSS.n1399 585
R856 VSS.n1398 VSS.n1397 585
R857 VSS.n1396 VSS.n1395 585
R858 VSS.n1394 VSS.n1393 585
R859 VSS.n1392 VSS.n1391 585
R860 VSS.n1390 VSS.n1389 585
R861 VSS.n1388 VSS.n1247 585
R862 VSS.n4784 VSS.n1247 585
R863 VSS.n1387 VSS.n1248 585
R864 VSS.n1508 VSS.n1507 585
R865 VSS.n1506 VSS.n1505 585
R866 VSS.n1504 VSS.n1503 585
R867 VSS.n1502 VSS.n1501 585
R868 VSS.n1500 VSS.n1499 585
R869 VSS.n1498 VSS.n1497 585
R870 VSS.n1496 VSS.n1495 585
R871 VSS.n1494 VSS.n1493 585
R872 VSS.n1492 VSS.n1491 585
R873 VSS.n1490 VSS.n1489 585
R874 VSS.n1511 VSS.n1510 585
R875 VSS.n1534 VSS.n1382 585
R876 VSS.n1533 VSS.n1532 585
R877 VSS.n1531 VSS.n1530 585
R878 VSS.n1529 VSS.n1528 585
R879 VSS.n1527 VSS.n1526 585
R880 VSS.n1525 VSS.n1524 585
R881 VSS.n1523 VSS.n1522 585
R882 VSS.n1521 VSS.n1520 585
R883 VSS.n1519 VSS.n1518 585
R884 VSS.n1517 VSS.n1516 585
R885 VSS.n1515 VSS.n1514 585
R886 VSS.n1513 VSS.n1512 585
R887 VSS.n1536 VSS.n1535 585
R888 VSS.n4788 VSS.n1219 585
R889 VSS.n4787 VSS.n4786 585
R890 VSS.n1221 VSS.n1220 585
R891 VSS.n1539 VSS.n1538 585
R892 VSS.n1541 VSS.n1540 585
R893 VSS.n1543 VSS.n1542 585
R894 VSS.n1545 VSS.n1544 585
R895 VSS.n1547 VSS.n1546 585
R896 VSS.n1549 VSS.n1548 585
R897 VSS.n1551 VSS.n1550 585
R898 VSS.n1553 VSS.n1552 585
R899 VSS.n1555 VSS.n1554 585
R900 VSS.n4788 VSS.n1218 585
R901 VSS.n4304 VSS.n4303 579.043
R902 VSS.n2620 VSS.n2588 578.947
R903 VSS.n2620 VSS.n2619 578.947
R904 VSS.n2619 VSS.n2618 578.947
R905 VSS.n2618 VSS.n2592 578.947
R906 VSS.n2592 VSS.n1742 578.947
R907 VSS.n2610 VSS.n1741 578.947
R908 VSS.n2610 VSS.n2609 578.947
R909 VSS.n2609 VSS.n2608 578.947
R910 VSS.n2608 VSS.n2597 578.947
R911 VSS.n2602 VSS.n2597 578.947
R912 VSS.n2602 VSS.n2601 578.947
R913 VSS.n2598 VSS.n2076 578.947
R914 VSS.n4016 VSS.n2076 578.947
R915 VSS.n4017 VSS.n4016 578.947
R916 VSS.n4019 VSS.n4017 578.947
R917 VSS.n4019 VSS.n4018 578.947
R918 VSS.n4026 VSS.n4025 578.947
R919 VSS.n4027 VSS.n4026 578.947
R920 VSS.n4027 VSS.n2069 578.947
R921 VSS.n4034 VSS.n2069 578.947
R922 VSS.n4035 VSS.n4034 578.947
R923 VSS.n4036 VSS.n4035 578.947
R924 VSS.n4038 VSS.n2063 578.947
R925 VSS.n4044 VSS.n2063 578.947
R926 VSS.n4045 VSS.n4044 578.947
R927 VSS.n4047 VSS.n4045 578.947
R928 VSS.n4047 VSS.n4046 578.947
R929 VSS.n4054 VSS.n4053 578.947
R930 VSS.n4056 VSS.n4054 578.947
R931 VSS.n4056 VSS.n4055 578.947
R932 VSS.n4055 VSS.n2056 578.947
R933 VSS.n4226 VSS.n2056 578.947
R934 VSS.n4227 VSS.n4226 578.947
R935 VSS.n4066 VSS.n4065 578.947
R936 VSS.n4218 VSS.n4066 578.947
R937 VSS.n4218 VSS.n4217 578.947
R938 VSS.n4217 VSS.n4216 578.947
R939 VSS.n4216 VSS.n4067 578.947
R940 VSS.n4210 VSS.n4209 578.947
R941 VSS.n4209 VSS.n4208 578.947
R942 VSS.n4208 VSS.n4071 578.947
R943 VSS.n4202 VSS.n4071 578.947
R944 VSS.n4202 VSS.n4201 578.947
R945 VSS.n4201 VSS.n4200 578.947
R946 VSS.n4082 VSS.n4081 578.947
R947 VSS.n4154 VSS.n4082 578.947
R948 VSS.n4154 VSS.n4153 578.947
R949 VSS.n4153 VSS.n4152 578.947
R950 VSS.n4152 VSS.n4083 578.947
R951 VSS.n4146 VSS.n4145 578.947
R952 VSS.n4145 VSS.n4144 578.947
R953 VSS.n4144 VSS.n4087 578.947
R954 VSS.n4138 VSS.n4087 578.947
R955 VSS.n4138 VSS.n4137 578.947
R956 VSS.n4137 VSS.n4136 578.947
R957 VSS.n4129 VSS.n4099 578.947
R958 VSS.n4129 VSS.n4128 578.947
R959 VSS.n4128 VSS.n4127 578.947
R960 VSS.n4127 VSS.n4100 578.947
R961 VSS.n4121 VSS.n4100 578.947
R962 VSS.n4119 VSS.n4118 578.947
R963 VSS.n4118 VSS.n4117 578.947
R964 VSS.n4117 VSS.n4105 578.947
R965 VSS.n4111 VSS.n4105 578.947
R966 VSS.n4111 VSS.n4110 578.947
R967 VSS.n4314 VSS.n4313 537.919
R968 VSS.n4296 VSS.t70 536.422
R969 VSS.n4329 VSS.n1746 530.74
R970 VSS.n4314 VSS.n4230 523.784
R971 VSS.t35 VSS.n1737 502.363
R972 VSS.n3175 VSS.t32 502.363
R973 VSS.n4638 VSS.t35 496.498
R974 VSS.n4672 VSS.t32 496.498
R975 VSS.n2601 VSS.n1702 482.457
R976 VSS.n4036 VSS.t32 482.457
R977 VSS.n4200 VSS.n4075 482.457
R978 VSS.n4136 VSS.n4091 482.457
R979 VSS.n4319 VSS.n1746 471.144
R980 VSS.n4282 VSS.n4281 454.401
R981 VSS.n4266 VSS.n4251 454.401
R982 VSS.n4256 VSS.n1245 434.791
R983 VSS.n4312 VSS.t70 406.812
R984 VSS.n2627 VSS.n2626 396.795
R985 VSS.n3121 VSS.n2627 396.795
R986 VSS.n3121 VSS.n3120 396.795
R987 VSS.n3120 VSS.n3119 396.795
R988 VSS.n3119 VSS.n2628 396.795
R989 VSS.n3110 VSS.n3109 396.795
R990 VSS.n3109 VSS.n3108 396.795
R991 VSS.n3108 VSS.n2637 396.795
R992 VSS.n3099 VSS.n2637 396.795
R993 VSS.n3099 VSS.n3098 396.795
R994 VSS.n3096 VSS.n2662 396.795
R995 VSS.n3086 VSS.n2662 396.795
R996 VSS.n3086 VSS.n3085 396.795
R997 VSS.n3085 VSS.n3084 396.795
R998 VSS.n3084 VSS.n2715 396.795
R999 VSS.n3075 VSS.n3074 396.795
R1000 VSS.n3074 VSS.n3073 396.795
R1001 VSS.n3073 VSS.n2724 396.795
R1002 VSS.n3064 VSS.n2724 396.795
R1003 VSS.n3064 VSS.n1740 396.795
R1004 VSS.n3055 VSS.n1739 396.795
R1005 VSS.n3055 VSS.n3054 396.795
R1006 VSS.n3054 VSS.n3053 396.795
R1007 VSS.n3053 VSS.n2782 396.795
R1008 VSS.n2802 VSS.n2782 396.795
R1009 VSS.n3040 VSS.n3039 396.795
R1010 VSS.n3039 VSS.n3038 396.795
R1011 VSS.n3038 VSS.n2803 396.795
R1012 VSS.n3029 VSS.n2803 396.795
R1013 VSS.n3029 VSS.n1753 396.795
R1014 VSS.n4637 VSS.n1754 396.795
R1015 VSS.n4466 VSS.n1754 396.795
R1016 VSS.n4467 VSS.n4466 396.795
R1017 VSS.n4469 VSS.n4467 396.795
R1018 VSS.n4469 VSS.n4468 396.795
R1019 VSS.n4484 VSS.n4456 396.795
R1020 VSS.n4485 VSS.n4484 396.795
R1021 VSS.n4487 VSS.n4485 396.795
R1022 VSS.n4487 VSS.n4486 396.795
R1023 VSS.n4486 VSS.n1750 396.795
R1024 VSS.n4363 VSS.n1751 396.795
R1025 VSS.n4363 VSS.n4362 396.795
R1026 VSS.n4362 VSS.n4361 396.795
R1027 VSS.n4361 VSS.n2003 396.795
R1028 VSS.n2028 VSS.n2003 396.795
R1029 VSS.n4348 VSS.n4347 396.795
R1030 VSS.n4347 VSS.n4346 396.795
R1031 VSS.n4346 VSS.n2029 396.795
R1032 VSS.n4337 VSS.n2029 396.795
R1033 VSS.n4337 VSS.n4336 396.795
R1034 VSS.n4303 VSS.t25 393.026
R1035 VSS.t35 VSS.n1742 392.399
R1036 VSS.n4018 VSS.t32 392.399
R1037 VSS.n4046 VSS.t32 392.399
R1038 VSS.n4067 VSS.t32 392.399
R1039 VSS.n4083 VSS.t32 392.399
R1040 VSS.n4121 VSS.t32 392.399
R1041 VSS.n4265 VSS.n4253 326.163
R1042 VSS.n4262 VSS.n4261 325.788
R1043 VSS.t25 VSS.n4302 316.322
R1044 VSS.n4274 VSS.n4252 311.416
R1045 VSS.n5354 VSS.n194 292.5
R1046 VSS.n5347 VSS.n5346 292.5
R1047 VSS.n5349 VSS.n203 292.5
R1048 VSS.n214 VSS.n202 292.5
R1049 VSS.n216 VSS.n215 292.5
R1050 VSS.n213 VSS.n206 292.5
R1051 VSS.n212 VSS.n211 292.5
R1052 VSS.n210 VSS.n209 292.5
R1053 VSS.n208 VSS.n207 292.5
R1054 VSS.n197 VSS.n195 292.5
R1055 VSS.n5353 VSS.n5352 292.5
R1056 VSS.n5345 VSS.n5344 292.5
R1057 VSS.n3648 VSS.n3642 292.5
R1058 VSS.n3650 VSS.n3641 292.5
R1059 VSS.n3653 VSS.n3652 292.5
R1060 VSS.n3655 VSS.n3654 292.5
R1061 VSS.n3657 VSS.n3639 292.5
R1062 VSS.n3659 VSS.n3638 292.5
R1063 VSS.n3662 VSS.n3661 292.5
R1064 VSS.n3664 VSS.n3663 292.5
R1065 VSS.n3666 VSS.n3632 292.5
R1066 VSS.n3669 VSS.n3668 292.5
R1067 VSS.n3670 VSS.n220 292.5
R1068 VSS.n5000 VSS.n4999 292.5
R1069 VSS.n4998 VSS.n4997 292.5
R1070 VSS.n4979 VSS.n4978 292.5
R1071 VSS.n4985 VSS.n4984 292.5
R1072 VSS.n4987 VSS.n4986 292.5
R1073 VSS.n4989 VSS.n4988 292.5
R1074 VSS.n4991 VSS.n4990 292.5
R1075 VSS.n4993 VSS.n4992 292.5
R1076 VSS.n4983 VSS.n4982 292.5
R1077 VSS.n4970 VSS.n4967 292.5
R1078 VSS.n5007 VSS.n5006 292.5
R1079 VSS.n5012 VSS.n699 292.5
R1080 VSS.n5014 VSS.n5013 292.5
R1081 VSS.n717 VSS.n716 292.5
R1082 VSS.n715 VSS.n714 292.5
R1083 VSS.n713 VSS.n712 292.5
R1084 VSS.n711 VSS.n710 292.5
R1085 VSS.n5017 VSS.n707 292.5
R1086 VSS.n5020 VSS.n5019 292.5
R1087 VSS.n5022 VSS.n5021 292.5
R1088 VSS.n5024 VSS.n5023 292.5
R1089 VSS.n705 VSS.n696 292.5
R1090 VSS.n5028 VSS.n5027 292.5
R1091 VSS.n4197 VSS.n4192 292.5
R1092 VSS.n1384 VSS.n1320 292.5
R1093 VSS.n1591 VSS.n1590 292.5
R1094 VSS.n1593 VSS.n1314 292.5
R1095 VSS.n1596 VSS.n1595 292.5
R1096 VSS.n1312 VSS.n1311 292.5
R1097 VSS.n1606 VSS.n1605 292.5
R1098 VSS.n1608 VSS.n1301 292.5
R1099 VSS.n1611 VSS.n1610 292.5
R1100 VSS.n1299 VSS.n1298 292.5
R1101 VSS.n4837 VSS.n4836 292.5
R1102 VSS.n1152 VSS.n1151 292.5
R1103 VSS.n1148 VSS.n1147 292.5
R1104 VSS.n1142 VSS.n1141 292.5
R1105 VSS.n1139 VSS.n1138 292.5
R1106 VSS.n1133 VSS.n1132 292.5
R1107 VSS.n1130 VSS.n761 292.5
R1108 VSS.n4924 VSS.n4923 292.5
R1109 VSS.n4927 VSS.n4926 292.5
R1110 VSS.n756 VSS.n748 292.5
R1111 VSS.n754 VSS.n747 292.5
R1112 VSS.n3566 VSS.n3565 292.5
R1113 VSS.n3562 VSS.n3561 292.5
R1114 VSS.n3542 VSS.n2316 292.5
R1115 VSS.n3544 VSS.n2315 292.5
R1116 VSS.n3547 VSS.n3546 292.5
R1117 VSS.n3540 VSS.n3539 292.5
R1118 VSS.n3874 VSS.n3873 292.5
R1119 VSS.n3876 VSS.n2261 292.5
R1120 VSS.n3879 VSS.n3878 292.5
R1121 VSS.n2267 VSS.n2266 292.5
R1122 VSS.n3780 VSS.n3779 292.5
R1123 VSS.n3776 VSS.n3775 292.5
R1124 VSS.n3770 VSS.n3769 292.5
R1125 VSS.n3767 VSS.n3766 292.5
R1126 VSS.n3761 VSS.n3760 292.5
R1127 VSS.n3758 VSS.n376 292.5
R1128 VSS.n5152 VSS.n5151 292.5
R1129 VSS.n5155 VSS.n5154 292.5
R1130 VSS.n568 VSS.n366 292.5
R1131 VSS.n570 VSS.n365 292.5
R1132 VSS.n566 VSS.n565 292.5
R1133 VSS.n562 VSS.n561 292.5
R1134 VSS.n551 VSS.n550 292.5
R1135 VSS.n548 VSS.n78 292.5
R1136 VSS.n546 VSS.n545 292.5
R1137 VSS.n5445 VSS.n5444 292.5
R1138 VSS.n5447 VSS.n70 292.5
R1139 VSS.n5450 VSS.n5449 292.5
R1140 VSS.n4193 VSS.n63 292.5
R1141 VSS.n4195 VSS.n62 292.5
R1142 VSS.n996 VSS.n959 292.5
R1143 VSS.n982 VSS.n981 292.5
R1144 VSS.n984 VSS.n983 292.5
R1145 VSS.n980 VSS.n971 292.5
R1146 VSS.n979 VSS.n978 292.5
R1147 VSS.n977 VSS.n976 292.5
R1148 VSS.n975 VSS.n974 292.5
R1149 VSS.n973 VSS.n972 292.5
R1150 VSS.n987 VSS.n968 292.5
R1151 VSS.n990 VSS.n989 292.5
R1152 VSS.n992 VSS.n991 292.5
R1153 VSS.n994 VSS.n993 292.5
R1154 VSS.n1011 VSS.n1010 292.5
R1155 VSS.n1013 VSS.n1005 292.5
R1156 VSS.n1016 VSS.n1015 292.5
R1157 VSS.n1018 VSS.n1017 292.5
R1158 VSS.n1020 VSS.n1003 292.5
R1159 VSS.n1022 VSS.n1002 292.5
R1160 VSS.n1025 VSS.n1024 292.5
R1161 VSS.n1027 VSS.n1026 292.5
R1162 VSS.n1029 VSS.n1000 292.5
R1163 VSS.n1031 VSS.n956 292.5
R1164 VSS.n1034 VSS.n1033 292.5
R1165 VSS.n1560 VSS.n1559 292.5
R1166 VSS.n1379 VSS.n1378 292.5
R1167 VSS.n1373 VSS.n1372 292.5
R1168 VSS.n1370 VSS.n1369 292.5
R1169 VSS.n1364 VSS.n1363 292.5
R1170 VSS.n1361 VSS.n1360 292.5
R1171 VSS.n1355 VSS.n1354 292.5
R1172 VSS.n4826 VSS.n4825 292.5
R1173 VSS.n4829 VSS.n4828 292.5
R1174 VSS.n1182 VSS.n1181 292.5
R1175 VSS.n1175 VSS.n1174 292.5
R1176 VSS.n1083 VSS.n1082 292.5
R1177 VSS.n1080 VSS.n1079 292.5
R1178 VSS.n1060 VSS.n1041 292.5
R1179 VSS.n1063 VSS.n1062 292.5
R1180 VSS.n1058 VSS.n1045 292.5
R1181 VSS.n1056 VSS.n1055 292.5
R1182 VSS.n1048 VSS.n1047 292.5
R1183 VSS.n4963 VSS.n4962 292.5
R1184 VSS.n4965 VSS.n720 292.5
R1185 VSS.n2302 VSS.n2301 292.5
R1186 VSS.n2298 VSS.n2297 292.5
R1187 VSS.n3616 VSS.n3615 292.5
R1188 VSS.n3619 VSS.n3618 292.5
R1189 VSS.n2291 VSS.n2290 292.5
R1190 VSS.n2288 VSS.n2284 292.5
R1191 VSS.n3839 VSS.n3838 292.5
R1192 VSS.n3841 VSS.n2279 292.5
R1193 VSS.n3844 VSS.n3843 292.5
R1194 VSS.n3810 VSS.n3809 292.5
R1195 VSS.n3803 VSS.n3802 292.5
R1196 VSS.n3699 VSS.n3672 292.5
R1197 VSS.n3702 VSS.n3701 292.5
R1198 VSS.n3697 VSS.n3675 292.5
R1199 VSS.n3695 VSS.n3694 292.5
R1200 VSS.n3682 VSS.n3681 292.5
R1201 VSS.n3679 VSS.n343 292.5
R1202 VSS.n3677 VSS.n342 292.5
R1203 VSS.n5172 VSS.n5171 292.5
R1204 VSS.n5175 VSS.n5174 292.5
R1205 VSS.n523 VSS.n522 292.5
R1206 VSS.n519 VSS.n518 292.5
R1207 VSS.n470 VSS.n469 292.5
R1208 VSS.n467 VSS.n39 292.5
R1209 VSS.n465 VSS.n464 292.5
R1210 VSS.n5466 VSS.n5465 292.5
R1211 VSS.n5468 VSS.n28 292.5
R1212 VSS.n5471 VSS.n5470 292.5
R1213 VSS.n4093 VSS.n21 292.5
R1214 VSS.n4095 VSS.n20 292.5
R1215 VSS.n4132 VSS.n4097 292.5
R1216 VSS.n266 VSS.n265 292.5
R1217 VSS.n264 VSS.n263 292.5
R1218 VSS.n245 VSS.n244 292.5
R1219 VSS.n251 VSS.n250 292.5
R1220 VSS.n253 VSS.n252 292.5
R1221 VSS.n255 VSS.n254 292.5
R1222 VSS.n257 VSS.n256 292.5
R1223 VSS.n259 VSS.n258 292.5
R1224 VSS.n249 VSS.n248 292.5
R1225 VSS.n575 VSS.n230 292.5
R1226 VSS.n235 VSS.n233 292.5
R1227 VSS.n5335 VSS.n5334 292.5
R1228 VSS.n595 VSS.n594 292.5
R1229 VSS.n593 VSS.n592 292.5
R1230 VSS.n591 VSS.n590 292.5
R1231 VSS.n589 VSS.n588 292.5
R1232 VSS.n587 VSS.n586 292.5
R1233 VSS.n598 VSS.n583 292.5
R1234 VSS.n601 VSS.n600 292.5
R1235 VSS.n603 VSS.n602 292.5
R1236 VSS.n605 VSS.n604 292.5
R1237 VSS.n581 VSS.n573 292.5
R1238 VSS.n609 VSS.n608 292.5
R1239 VSS.n5363 VSS.n163 292.5
R1240 VSS.n5365 VSS.n5364 292.5
R1241 VSS.n179 VSS.n178 292.5
R1242 VSS.n177 VSS.n176 292.5
R1243 VSS.n175 VSS.n174 292.5
R1244 VSS.n173 VSS.n172 292.5
R1245 VSS.n5368 VSS.n169 292.5
R1246 VSS.n5371 VSS.n5370 292.5
R1247 VSS.n5373 VSS.n5372 292.5
R1248 VSS.n5375 VSS.n5374 292.5
R1249 VSS.n5033 VSS.n676 292.5
R1250 VSS.n5035 VSS.n5034 292.5
R1251 VSS.n692 VSS.n691 292.5
R1252 VSS.n690 VSS.n689 292.5
R1253 VSS.n688 VSS.n687 292.5
R1254 VSS.n686 VSS.n685 292.5
R1255 VSS.n5038 VSS.n682 292.5
R1256 VSS.n5041 VSS.n5040 292.5
R1257 VSS.n5043 VSS.n5042 292.5
R1258 VSS.n5045 VSS.n5044 292.5
R1259 VSS.n4842 VSS.n869 292.5
R1260 VSS.n4844 VSS.n4843 292.5
R1261 VSS.n885 VSS.n884 292.5
R1262 VSS.n883 VSS.n882 292.5
R1263 VSS.n881 VSS.n880 292.5
R1264 VSS.n879 VSS.n878 292.5
R1265 VSS.n4847 VSS.n875 292.5
R1266 VSS.n4850 VSS.n4849 292.5
R1267 VSS.n4852 VSS.n4851 292.5
R1268 VSS.n4854 VSS.n4853 292.5
R1269 VSS.n3169 VSS.n3164 292.5
R1270 VSS.n3165 VSS.n3164 292.5
R1271 VSS.n3170 VSS.n3162 292.5
R1272 VSS.n3162 VSS.n3161 292.5
R1273 VSS.n3172 VSS.n3171 292.5
R1274 VSS.n3173 VSS.n3172 292.5
R1275 VSS.n3163 VSS.n3159 292.5
R1276 VSS.n3174 VSS.n3159 292.5
R1277 VSS.n3176 VSS.n3160 292.5
R1278 VSS.n3176 VSS.n3175 292.5
R1279 VSS.n3177 VSS.n3158 292.5
R1280 VSS.n3178 VSS.n3177 292.5
R1281 VSS.n3181 VSS.n3180 292.5
R1282 VSS.n3180 VSS.n3179 292.5
R1283 VSS.n3182 VSS.n3157 292.5
R1284 VSS.n3157 VSS.n3156 292.5
R1285 VSS.n3184 VSS.n3183 292.5
R1286 VSS.n3185 VSS.n3184 292.5
R1287 VSS.n3168 VSS.n3167 292.5
R1288 VSS.n3167 VSS.n3166 292.5
R1289 VSS.n2203 VSS.n2202 292.5
R1290 VSS.n2201 VSS.n2178 292.5
R1291 VSS.n2200 VSS.n2199 292.5
R1292 VSS.n2181 VSS.n2180 292.5
R1293 VSS.n2189 VSS.n2188 292.5
R1294 VSS.n2191 VSS.n2190 292.5
R1295 VSS.n2193 VSS.n2192 292.5
R1296 VSS.n2195 VSS.n2194 292.5
R1297 VSS.n2187 VSS.n2184 292.5
R1298 VSS.n2186 VSS.n2185 292.5
R1299 VSS.n2206 VSS.n2172 292.5
R1300 VSS.n3411 VSS.n3393 292.5
R1301 VSS.n3413 VSS.n3412 292.5
R1302 VSS.n3410 VSS.n3397 292.5
R1303 VSS.n3409 VSS.n3408 292.5
R1304 VSS.n3407 VSS.n3406 292.5
R1305 VSS.n3405 VSS.n3404 292.5
R1306 VSS.n3403 VSS.n3402 292.5
R1307 VSS.n3401 VSS.n3400 292.5
R1308 VSS.n3399 VSS.n3398 292.5
R1309 VSS.n3417 VSS.n2216 292.5
R1310 VSS.n3932 VSS.n3930 292.5
R1311 VSS.n3934 VSS.n3929 292.5
R1312 VSS.n3937 VSS.n3936 292.5
R1313 VSS.n3939 VSS.n3938 292.5
R1314 VSS.n3941 VSS.n3927 292.5
R1315 VSS.n3943 VSS.n3926 292.5
R1316 VSS.n3946 VSS.n3945 292.5
R1317 VSS.n3948 VSS.n3947 292.5
R1318 VSS.n3950 VSS.n3924 292.5
R1319 VSS.n3952 VSS.n3921 292.5
R1320 VSS.n3955 VSS.n3954 292.5
R1321 VSS.n5054 VSS.n191 292.5
R1322 VSS.n5072 VSS.n5071 292.5
R1323 VSS.n5070 VSS.n5069 292.5
R1324 VSS.n5068 VSS.n5067 292.5
R1325 VSS.n5066 VSS.n5065 292.5
R1326 VSS.n5064 VSS.n5063 292.5
R1327 VSS.n5075 VSS.n5060 292.5
R1328 VSS.n5078 VSS.n5077 292.5
R1329 VSS.n5080 VSS.n5079 292.5
R1330 VSS.n5082 VSS.n5081 292.5
R1331 VSS.n4557 VSS.n4556 292.5
R1332 VSS.n4555 VSS.n4534 292.5
R1333 VSS.n4554 VSS.n4553 292.5
R1334 VSS.n4537 VSS.n4536 292.5
R1335 VSS.n4543 VSS.n4542 292.5
R1336 VSS.n4545 VSS.n4544 292.5
R1337 VSS.n4547 VSS.n4546 292.5
R1338 VSS.n4549 VSS.n4548 292.5
R1339 VSS.n4541 VSS.n4540 292.5
R1340 VSS.n4529 VSS.n1951 292.5
R1341 VSS.n4561 VSS.n4560 292.5
R1342 VSS.n2984 VSS.n2965 292.5
R1343 VSS.n2986 VSS.n2985 292.5
R1344 VSS.n2982 VSS.n2981 292.5
R1345 VSS.n2980 VSS.n2979 292.5
R1346 VSS.n2978 VSS.n2977 292.5
R1347 VSS.n2976 VSS.n2975 292.5
R1348 VSS.n2989 VSS.n2972 292.5
R1349 VSS.n2992 VSS.n2991 292.5
R1350 VSS.n2994 VSS.n2993 292.5
R1351 VSS.n2996 VSS.n2995 292.5
R1352 VSS.n2941 VSS.n2940 292.5
R1353 VSS.n2943 VSS.n2942 292.5
R1354 VSS.n2945 VSS.n2937 292.5
R1355 VSS.n2947 VSS.n2936 292.5
R1356 VSS.n2950 VSS.n2949 292.5
R1357 VSS.n2952 VSS.n2951 292.5
R1358 VSS.n2954 VSS.n2934 292.5
R1359 VSS.n2956 VSS.n2933 292.5
R1360 VSS.n2959 VSS.n2958 292.5
R1361 VSS.n2961 VSS.n2960 292.5
R1362 VSS.n2963 VSS.n2330 292.5
R1363 VSS.n4566 VSS.n4565 292.5
R1364 VSS.n1887 VSS.n1864 292.5
R1365 VSS.n4574 VSS.n4573 292.5
R1366 VSS.n4577 VSS.n4576 292.5
R1367 VSS.n1860 VSS.n1859 292.5
R1368 VSS.n1857 VSS.n1851 292.5
R1369 VSS.n4591 VSS.n4590 292.5
R1370 VSS.n4593 VSS.n1843 292.5
R1371 VSS.n4596 VSS.n4595 292.5
R1372 VSS.n2327 VSS.n2326 292.5
R1373 VSS.n3441 VSS.n2323 292.5
R1374 VSS.n3439 VSS.n3438 292.5
R1375 VSS.n2375 VSS.n2374 292.5
R1376 VSS.n2372 VSS.n2371 292.5
R1377 VSS.n2366 VSS.n2365 292.5
R1378 VSS.n2363 VSS.n2362 292.5
R1379 VSS.n2357 VSS.n2356 292.5
R1380 VSS.n2354 VSS.n2353 292.5
R1381 VSS.n3917 VSS.n3916 292.5
R1382 VSS.n3919 VSS.n2218 292.5
R1383 VSS.n3313 VSS.n3312 292.5
R1384 VSS.n3309 VSS.n3228 292.5
R1385 VSS.n3321 VSS.n3320 292.5
R1386 VSS.n3324 VSS.n3323 292.5
R1387 VSS.n3224 VSS.n3223 292.5
R1388 VSS.n3221 VSS.n3215 292.5
R1389 VSS.n3338 VSS.n3337 292.5
R1390 VSS.n3340 VSS.n3208 292.5
R1391 VSS.n3343 VSS.n3342 292.5
R1392 VSS.n3205 VSS.n3204 292.5
R1393 VSS.n3968 VSS.n3967 292.5
R1394 VSS.n3970 VSS.n2145 292.5
R1395 VSS.n3973 VSS.n3972 292.5
R1396 VSS.n2142 VSS.n2139 292.5
R1397 VSS.n3981 VSS.n3980 292.5
R1398 VSS.n3984 VSS.n3983 292.5
R1399 VSS.n2132 VSS.n2125 292.5
R1400 VSS.n2130 VSS.n2124 292.5
R1401 VSS.n3994 VSS.n3993 292.5
R1402 VSS.n3997 VSS.n3996 292.5
R1403 VSS.n2757 VSS.n2755 292.5
R1404 VSS.n2760 VSS.n2759 292.5
R1405 VSS.n2762 VSS.n2761 292.5
R1406 VSS.n2764 VSS.n2753 292.5
R1407 VSS.n2766 VSS.n2752 292.5
R1408 VSS.n2769 VSS.n2768 292.5
R1409 VSS.n2771 VSS.n2770 292.5
R1410 VSS.n2773 VSS.n2749 292.5
R1411 VSS.n2776 VSS.n2775 292.5
R1412 VSS.n3003 VSS.n2817 292.5
R1413 VSS.n3006 VSS.n3005 292.5
R1414 VSS.n3008 VSS.n3007 292.5
R1415 VSS.n3010 VSS.n2815 292.5
R1416 VSS.n3012 VSS.n2814 292.5
R1417 VSS.n3015 VSS.n3014 292.5
R1418 VSS.n3017 VSS.n3016 292.5
R1419 VSS.n3019 VSS.n2811 292.5
R1420 VSS.n3022 VSS.n3021 292.5
R1421 VSS.n4519 VSS.n4518 292.5
R1422 VSS.n4517 VSS.n4516 292.5
R1423 VSS.n4514 VSS.n1992 292.5
R1424 VSS.n4512 VSS.n4511 292.5
R1425 VSS.n4510 VSS.n4509 292.5
R1426 VSS.n4507 VSS.n1994 292.5
R1427 VSS.n4505 VSS.n4504 292.5
R1428 VSS.n4503 VSS.n4502 292.5
R1429 VSS.n4500 VSS.n1996 292.5
R1430 VSS.n4526 VSS.n1955 292.5
R1431 VSS.n1980 VSS.n1979 292.5
R1432 VSS.n1982 VSS.n1981 292.5
R1433 VSS.n1978 VSS.n1969 292.5
R1434 VSS.n1977 VSS.n1976 292.5
R1435 VSS.n1975 VSS.n1974 292.5
R1436 VSS.n1973 VSS.n1972 292.5
R1437 VSS.n1971 VSS.n1970 292.5
R1438 VSS.n1985 VSS.n1966 292.5
R1439 VSS.n1988 VSS.n1987 292.5
R1440 VSS.n2676 VSS.n2674 292.5
R1441 VSS.n2674 VSS.n2673 292.5
R1442 VSS.n2678 VSS.n2677 292.5
R1443 VSS.n2679 VSS.n2678 292.5
R1444 VSS.n2675 VSS.n2671 292.5
R1445 VSS.n2680 VSS.n2671 292.5
R1446 VSS.n2682 VSS.n2672 292.5
R1447 VSS.n2682 VSS.n2681 292.5
R1448 VSS.n2683 VSS.n2670 292.5
R1449 VSS.n2683 VSS.n1737 292.5
R1450 VSS.n2685 VSS.n2684 292.5
R1451 VSS.n2684 VSS.n1736 292.5
R1452 VSS.n2686 VSS.n2668 292.5
R1453 VSS.n2668 VSS.n2667 292.5
R1454 VSS.n2688 VSS.n2687 292.5
R1455 VSS.n2689 VSS.n2688 292.5
R1456 VSS.n2669 VSS.n2666 292.5
R1457 VSS.n2690 VSS.n2666 292.5
R1458 VSS.n2692 VSS.n2691 292.5
R1459 VSS.n2696 VSS.n2661 292.5
R1460 VSS.n2496 VSS.n1738 292.5
R1461 VSS.n4686 VSS.n4685 292.5
R1462 VSS.n1818 VSS.n1817 292.5
R1463 VSS.n1824 VSS.n1823 292.5
R1464 VSS.n1813 VSS.n1786 292.5
R1465 VSS.n1808 VSS.n1807 292.5
R1466 VSS.n1803 VSS.n1802 292.5
R1467 VSS.n1797 VSS.n1796 292.5
R1468 VSS.n1792 VSS.n1791 292.5
R1469 VSS.n1782 VSS.n1645 292.5
R1470 VSS.n1671 VSS.n1644 292.5
R1471 VSS.n4690 VSS.n4689 292.5
R1472 VSS.n1677 VSS.n1667 292.5
R1473 VSS.n4433 VSS.n1706 292.5
R1474 VSS.n4432 VSS.n4431 292.5
R1475 VSS.n4425 VSS.n4424 292.5
R1476 VSS.n4422 VSS.n4421 292.5
R1477 VSS.n4416 VSS.n4415 292.5
R1478 VSS.n4413 VSS.n4412 292.5
R1479 VSS.n4407 VSS.n4406 292.5
R1480 VSS.n4404 VSS.n4403 292.5
R1481 VSS.n4623 VSS.n4622 292.5
R1482 VSS.n4626 VSS.n4625 292.5
R1483 VSS.n2925 VSS.n2924 292.5
R1484 VSS.n2927 VSS.n1683 292.5
R1485 VSS.n2902 VSS.n1705 292.5
R1486 VSS.n2900 VSS.n2899 292.5
R1487 VSS.n2893 VSS.n2892 292.5
R1488 VSS.n2890 VSS.n2889 292.5
R1489 VSS.n2884 VSS.n2883 292.5
R1490 VSS.n2881 VSS.n2880 292.5
R1491 VSS.n2875 VSS.n2874 292.5
R1492 VSS.n2872 VSS.n2871 292.5
R1493 VSS.n2866 VSS.n2865 292.5
R1494 VSS.n2863 VSS.n2396 292.5
R1495 VSS.n2395 VSS.n2394 292.5
R1496 VSS.n3421 VSS.n1689 292.5
R1497 VSS.n3384 VSS.n1704 292.5
R1498 VSS.n3382 VSS.n3381 292.5
R1499 VSS.n3266 VSS.n3265 292.5
R1500 VSS.n3263 VSS.n3262 292.5
R1501 VSS.n3257 VSS.n3256 292.5
R1502 VSS.n3254 VSS.n3253 292.5
R1503 VSS.n3248 VSS.n3247 292.5
R1504 VSS.n3245 VSS.n3244 292.5
R1505 VSS.n3370 VSS.n3369 292.5
R1506 VSS.n3373 VSS.n3372 292.5
R1507 VSS.n3192 VSS.n3191 292.5
R1508 VSS.n3189 VSS.n1695 292.5
R1509 VSS.n3152 VSS.n1703 292.5
R1510 VSS.n3150 VSS.n3149 292.5
R1511 VSS.n2558 VSS.n2557 292.5
R1512 VSS.n2561 VSS.n2560 292.5
R1513 VSS.n2551 VSS.n2550 292.5
R1514 VSS.n2548 VSS.n2547 292.5
R1515 VSS.n2571 VSS.n2570 292.5
R1516 VSS.n2574 VSS.n2573 292.5
R1517 VSS.n2539 VSS.n2538 292.5
R1518 VSS.n2536 VSS.n2535 292.5
R1519 VSS.n4009 VSS.n4008 292.5
R1520 VSS.n4011 VSS.n1701 292.5
R1521 VSS.n3186 VSS.n2495 292.5
R1522 VSS.n1916 VSS.n1254 292.5
R1523 VSS.n1919 VSS.n1918 292.5
R1524 VSS.n1928 VSS.n1927 292.5
R1525 VSS.n1930 VSS.n1905 292.5
R1526 VSS.n1933 VSS.n1932 292.5
R1527 VSS.n1903 VSS.n1902 292.5
R1528 VSS.n1942 VSS.n1941 292.5
R1529 VSS.n1944 VSS.n1892 292.5
R1530 VSS.n1946 VSS.n1622 292.5
R1531 VSS.n1948 VSS.n1621 292.5
R1532 VSS.n1484 VSS.n1407 292.5
R1533 VSS.n1482 VSS.n1481 292.5
R1534 VSS.n1425 VSS.n1410 292.5
R1535 VSS.n1427 VSS.n1411 292.5
R1536 VSS.n1429 VSS.n1412 292.5
R1537 VSS.n1432 VSS.n1431 292.5
R1538 VSS.n1423 VSS.n1422 292.5
R1539 VSS.n1417 VSS.n1416 292.5
R1540 VSS.n4768 VSS.n4767 292.5
R1541 VSS.n4771 VSS.n4770 292.5
R1542 VSS.n4742 VSS.n4741 292.5
R1543 VSS.n4739 VSS.n4738 292.5
R1544 VSS.n4860 VSS.n4859 292.5
R1545 VSS.n4863 VSS.n4862 292.5
R1546 VSS.n861 VSS.n856 292.5
R1547 VSS.n859 VSS.n855 292.5
R1548 VSS.n4873 VSS.n4872 292.5
R1549 VSS.n4876 VSS.n4875 292.5
R1550 VSS.n845 VSS.n841 292.5
R1551 VSS.n843 VSS.n840 292.5
R1552 VSS.n4886 VSS.n4885 292.5
R1553 VSS.n4888 VSS.n783 292.5
R1554 VSS.n4890 VSS.n782 292.5
R1555 VSS.n4893 VSS.n4892 292.5
R1556 VSS.n670 VSS.n668 292.5
R1557 VSS.n3510 VSS.n3509 292.5
R1558 VSS.n3506 VSS.n3505 292.5
R1559 VSS.n3486 VSS.n3467 292.5
R1560 VSS.n3489 VSS.n3488 292.5
R1561 VSS.n3484 VSS.n3483 292.5
R1562 VSS.n3478 VSS.n3477 292.5
R1563 VSS.n3475 VSS.n3474 292.5
R1564 VSS.n3906 VSS.n3905 292.5
R1565 VSS.n3909 VSS.n3908 292.5
R1566 VSS.n2422 VSS.n2421 292.5
R1567 VSS.n663 VSS.n662 292.5
R1568 VSS.n5088 VSS.n5087 292.5
R1569 VSS.n5091 VSS.n5090 292.5
R1570 VSS.n654 VSS.n649 292.5
R1571 VSS.n652 VSS.n648 292.5
R1572 VSS.n5101 VSS.n5100 292.5
R1573 VSS.n5104 VSS.n5103 292.5
R1574 VSS.n638 VSS.n634 292.5
R1575 VSS.n636 VSS.n633 292.5
R1576 VSS.n5114 VSS.n5113 292.5
R1577 VSS.n5116 VSS.n398 292.5
R1578 VSS.n5118 VSS.n397 292.5
R1579 VSS.n5121 VSS.n5120 292.5
R1580 VSS.n5381 VSS.n5380 292.5
R1581 VSS.n5384 VSS.n5383 292.5
R1582 VSS.n154 VSS.n149 292.5
R1583 VSS.n152 VSS.n148 292.5
R1584 VSS.n5394 VSS.n5393 292.5
R1585 VSS.n5397 VSS.n5396 292.5
R1586 VSS.n138 VSS.n134 292.5
R1587 VSS.n136 VSS.n133 292.5
R1588 VSS.n5407 VSS.n5406 292.5
R1589 VSS.n5409 VSS.n102 292.5
R1590 VSS.n5411 VSS.n101 292.5
R1591 VSS.n5414 VSS.n5413 292.5
R1592 VSS.n5329 VSS.n5328 292.5
R1593 VSS.n5329 VSS.n271 292.5
R1594 VSS.n5329 VSS.n270 292.5
R1595 VSS.n5330 VSS.n5329 292.5
R1596 VSS.n4267 VSS.n4248 292.5
R1597 VSS.t21 VSS.n4248 292.5
R1598 VSS.n4284 VSS.n4283 292.5
R1599 VSS.t21 VSS.n4284 292.5
R1600 VSS.n4299 VSS.t27 284.457
R1601 VSS.n4305 VSS.n4292 284.455
R1602 VSS.n4300 VSS.t37 284.216
R1603 VSS.n4784 VSS.n4783 277.688
R1604 VSS.n4784 VSS.n1227 277.688
R1605 VSS.n4784 VSS.n1239 277.688
R1606 VSS.n5348 VSS.n218 272.089
R1607 VSS.n5350 VSS.n201 272.089
R1608 VSS.n218 VSS.n217 272.089
R1609 VSS.n5350 VSS.n200 272.089
R1610 VSS.n218 VSS.n205 272.089
R1611 VSS.n5350 VSS.n199 272.089
R1612 VSS.n218 VSS.n204 272.089
R1613 VSS.n5351 VSS.n5350 272.089
R1614 VSS.n218 VSS.n196 272.089
R1615 VSS.n5350 VSS.n198 272.089
R1616 VSS.n3649 VSS.n3634 272.089
R1617 VSS.n3647 VSS.n3636 272.089
R1618 VSS.n3651 VSS.n3636 272.089
R1619 VSS.n3640 VSS.n3634 272.089
R1620 VSS.n3656 VSS.n3636 272.089
R1621 VSS.n3658 VSS.n3634 272.089
R1622 VSS.n3660 VSS.n3636 272.089
R1623 VSS.n3637 VSS.n3634 272.089
R1624 VSS.n3665 VSS.n3636 272.089
R1625 VSS.n3667 VSS.n3634 272.089
R1626 VSS.n3636 VSS.n3633 272.089
R1627 VSS.n4995 VSS.n4977 272.089
R1628 VSS.n5005 VSS.n4975 272.089
R1629 VSS.n4996 VSS.n4995 272.089
R1630 VSS.n5005 VSS.n4974 272.089
R1631 VSS.n4995 VSS.n4980 272.089
R1632 VSS.n5005 VSS.n4973 272.089
R1633 VSS.n4995 VSS.n4981 272.089
R1634 VSS.n5005 VSS.n4972 272.089
R1635 VSS.n4995 VSS.n4994 272.089
R1636 VSS.n5005 VSS.n4971 272.089
R1637 VSS.n4995 VSS.n4969 272.089
R1638 VSS.n5016 VSS.n5015 272.089
R1639 VSS.n5026 VSS.n701 272.089
R1640 VSS.n5016 VSS.n709 272.089
R1641 VSS.n5026 VSS.n702 272.089
R1642 VSS.n5016 VSS.n708 272.089
R1643 VSS.n5026 VSS.n703 272.089
R1644 VSS.n5018 VSS.n5016 272.089
R1645 VSS.n5026 VSS.n704 272.089
R1646 VSS.n5016 VSS.n706 272.089
R1647 VSS.n5026 VSS.n5025 272.089
R1648 VSS.n5016 VSS.n698 272.089
R1649 VSS.n4194 VSS.n69 272.089
R1650 VSS.n5448 VSS.n69 272.089
R1651 VSS.n72 VSS.n69 272.089
R1652 VSS.n549 VSS.n69 272.089
R1653 VSS.n563 VSS.n69 272.089
R1654 VSS.n571 VSS.n69 272.089
R1655 VSS.n372 VSS.n69 272.089
R1656 VSS.n373 VSS.n69 272.089
R1657 VSS.n3756 VSS.n69 272.089
R1658 VSS.n3752 VSS.n69 272.089
R1659 VSS.n3778 VSS.n69 272.089
R1660 VSS.n193 VSS.n69 272.089
R1661 VSS.n3877 VSS.n69 272.089
R1662 VSS.n2262 VSS.n69 272.089
R1663 VSS.n3545 VSS.n69 272.089
R1664 VSS.n2310 VSS.n69 272.089
R1665 VSS.n3564 VSS.n69 272.089
R1666 VSS.n695 VSS.n69 272.089
R1667 VSS.n757 VSS.n69 272.089
R1668 VSS.n758 VSS.n69 272.089
R1669 VSS.n1128 VSS.n69 272.089
R1670 VSS.n1124 VSS.n69 272.089
R1671 VSS.n1150 VSS.n69 272.089
R1672 VSS.n889 VSS.n69 272.089
R1673 VSS.n1609 VSS.n69 272.089
R1674 VSS.n1302 VSS.n69 272.089
R1675 VSS.n1594 VSS.n69 272.089
R1676 VSS.n1315 VSS.n69 272.089
R1677 VSS.n1385 VSS.n71 272.089
R1678 VSS.n1592 VSS.n71 272.089
R1679 VSS.n1313 VSS.n71 272.089
R1680 VSS.n1607 VSS.n71 272.089
R1681 VSS.n1300 VSS.n71 272.089
R1682 VSS.n4838 VSS.n71 272.089
R1683 VSS.n1149 VSS.n71 272.089
R1684 VSS.n1140 VSS.n71 272.089
R1685 VSS.n1131 VSS.n71 272.089
R1686 VSS.n4925 VSS.n71 272.089
R1687 VSS.n755 VSS.n71 272.089
R1688 VSS.n3563 VSS.n71 272.089
R1689 VSS.n3543 VSS.n71 272.089
R1690 VSS.n3541 VSS.n71 272.089
R1691 VSS.n3875 VSS.n71 272.089
R1692 VSS.n2259 VSS.n71 272.089
R1693 VSS.n3777 VSS.n71 272.089
R1694 VSS.n3768 VSS.n71 272.089
R1695 VSS.n3759 VSS.n71 272.089
R1696 VSS.n5153 VSS.n71 272.089
R1697 VSS.n569 VSS.n71 272.089
R1698 VSS.n564 VSS.n71 272.089
R1699 VSS.n544 VSS.n71 272.089
R1700 VSS.n547 VSS.n71 272.089
R1701 VSS.n5446 VSS.n71 272.089
R1702 VSS.n71 VSS.n68 272.089
R1703 VSS.n4196 VSS.n71 272.089
R1704 VSS.n986 VSS.n957 272.089
R1705 VSS.n995 VSS.n961 272.089
R1706 VSS.n986 VSS.n985 272.089
R1707 VSS.n995 VSS.n962 272.089
R1708 VSS.n986 VSS.n970 272.089
R1709 VSS.n995 VSS.n963 272.089
R1710 VSS.n986 VSS.n969 272.089
R1711 VSS.n995 VSS.n964 272.089
R1712 VSS.n988 VSS.n986 272.089
R1713 VSS.n995 VSS.n965 272.089
R1714 VSS.n986 VSS.n967 272.089
R1715 VSS.n1012 VSS.n998 272.089
R1716 VSS.n1007 VSS.n999 272.089
R1717 VSS.n1014 VSS.n999 272.089
R1718 VSS.n1004 VSS.n998 272.089
R1719 VSS.n1019 VSS.n999 272.089
R1720 VSS.n1021 VSS.n998 272.089
R1721 VSS.n1023 VSS.n999 272.089
R1722 VSS.n1001 VSS.n998 272.089
R1723 VSS.n1028 VSS.n999 272.089
R1724 VSS.n1030 VSS.n998 272.089
R1725 VSS.n1032 VSS.n999 272.089
R1726 VSS.n4094 VSS.n27 272.089
R1727 VSS.n5469 VSS.n27 272.089
R1728 VSS.n30 VSS.n27 272.089
R1729 VSS.n468 VSS.n27 272.089
R1730 VSS.n520 VSS.n27 272.089
R1731 VSS.n232 VSS.n27 272.089
R1732 VSS.n338 VSS.n27 272.089
R1733 VSS.n3680 VSS.n27 272.089
R1734 VSS.n3696 VSS.n27 272.089
R1735 VSS.n3700 VSS.n27 272.089
R1736 VSS.n3804 VSS.n27 272.089
R1737 VSS.n3808 VSS.n27 272.089
R1738 VSS.n3842 VSS.n27 272.089
R1739 VSS.n2280 VSS.n27 272.089
R1740 VSS.n2292 VSS.n27 272.089
R1741 VSS.n2293 VSS.n27 272.089
R1742 VSS.n2300 VSS.n27 272.089
R1743 VSS.n4966 VSS.n27 272.089
R1744 VSS.n721 VSS.n27 272.089
R1745 VSS.n1057 VSS.n27 272.089
R1746 VSS.n1061 VSS.n27 272.089
R1747 VSS.n1081 VSS.n27 272.089
R1748 VSS.n1176 VSS.n27 272.089
R1749 VSS.n914 VSS.n27 272.089
R1750 VSS.n915 VSS.n27 272.089
R1751 VSS.n1362 VSS.n27 272.089
R1752 VSS.n1371 VSS.n27 272.089
R1753 VSS.n1380 VSS.n27 272.089
R1754 VSS.n1558 VSS.n29 272.089
R1755 VSS.n1343 VSS.n29 272.089
R1756 VSS.n1347 VSS.n29 272.089
R1757 VSS.n1353 VSS.n29 272.089
R1758 VSS.n4827 VSS.n29 272.089
R1759 VSS.n1180 VSS.n29 272.089
R1760 VSS.n1035 VSS.n29 272.089
R1761 VSS.n1040 VSS.n29 272.089
R1762 VSS.n1059 VSS.n29 272.089
R1763 VSS.n1046 VSS.n29 272.089
R1764 VSS.n4964 VSS.n29 272.089
R1765 VSS.n2299 VSS.n29 272.089
R1766 VSS.n3617 VSS.n29 272.089
R1767 VSS.n2289 VSS.n29 272.089
R1768 VSS.n3840 VSS.n29 272.089
R1769 VSS.n2277 VSS.n29 272.089
R1770 VSS.n3671 VSS.n29 272.089
R1771 VSS.n3698 VSS.n29 272.089
R1772 VSS.n3676 VSS.n29 272.089
R1773 VSS.n3678 VSS.n29 272.089
R1774 VSS.n5173 VSS.n29 272.089
R1775 VSS.n521 VSS.n29 272.089
R1776 VSS.n460 VSS.n29 272.089
R1777 VSS.n466 VSS.n29 272.089
R1778 VSS.n5467 VSS.n29 272.089
R1779 VSS.n29 VSS.n26 272.089
R1780 VSS.n4096 VSS.n29 272.089
R1781 VSS.n261 VSS.n242 272.089
R1782 VSS.n5333 VSS.n240 272.089
R1783 VSS.n262 VSS.n261 272.089
R1784 VSS.n5333 VSS.n239 272.089
R1785 VSS.n261 VSS.n246 272.089
R1786 VSS.n5333 VSS.n238 272.089
R1787 VSS.n261 VSS.n247 272.089
R1788 VSS.n5333 VSS.n237 272.089
R1789 VSS.n261 VSS.n260 272.089
R1790 VSS.n5333 VSS.n236 272.089
R1791 VSS.n597 VSS.n596 272.089
R1792 VSS.n261 VSS.n234 272.089
R1793 VSS.n607 VSS.n577 272.089
R1794 VSS.n597 VSS.n585 272.089
R1795 VSS.n607 VSS.n578 272.089
R1796 VSS.n597 VSS.n584 272.089
R1797 VSS.n607 VSS.n579 272.089
R1798 VSS.n599 VSS.n597 272.089
R1799 VSS.n607 VSS.n580 272.089
R1800 VSS.n597 VSS.n582 272.089
R1801 VSS.n607 VSS.n606 272.089
R1802 VSS.n597 VSS.n574 272.089
R1803 VSS.n5367 VSS.n5366 272.089
R1804 VSS.n5377 VSS.n164 272.089
R1805 VSS.n5367 VSS.n171 272.089
R1806 VSS.n5377 VSS.n165 272.089
R1807 VSS.n5367 VSS.n170 272.089
R1808 VSS.n5377 VSS.n166 272.089
R1809 VSS.n5369 VSS.n5367 272.089
R1810 VSS.n5377 VSS.n167 272.089
R1811 VSS.n5367 VSS.n168 272.089
R1812 VSS.n5377 VSS.n5376 272.089
R1813 VSS.n5037 VSS.n5036 272.089
R1814 VSS.n5047 VSS.n677 272.089
R1815 VSS.n5037 VSS.n684 272.089
R1816 VSS.n5047 VSS.n678 272.089
R1817 VSS.n5037 VSS.n683 272.089
R1818 VSS.n5047 VSS.n679 272.089
R1819 VSS.n5039 VSS.n5037 272.089
R1820 VSS.n5047 VSS.n680 272.089
R1821 VSS.n5037 VSS.n681 272.089
R1822 VSS.n5047 VSS.n5046 272.089
R1823 VSS.n4846 VSS.n4845 272.089
R1824 VSS.n4856 VSS.n870 272.089
R1825 VSS.n4846 VSS.n877 272.089
R1826 VSS.n4856 VSS.n871 272.089
R1827 VSS.n4846 VSS.n876 272.089
R1828 VSS.n4856 VSS.n872 272.089
R1829 VSS.n4848 VSS.n4846 272.089
R1830 VSS.n4856 VSS.n873 272.089
R1831 VSS.n4846 VSS.n874 272.089
R1832 VSS.n4856 VSS.n4855 272.089
R1833 VSS.n2197 VSS.n2179 272.089
R1834 VSS.n2205 VSS.n2204 272.089
R1835 VSS.n2198 VSS.n2197 272.089
R1836 VSS.n2205 VSS.n2177 272.089
R1837 VSS.n2197 VSS.n2182 272.089
R1838 VSS.n2205 VSS.n2176 272.089
R1839 VSS.n2197 VSS.n2183 272.089
R1840 VSS.n2205 VSS.n2175 272.089
R1841 VSS.n2197 VSS.n2196 272.089
R1842 VSS.n2205 VSS.n2174 272.089
R1843 VSS.n2197 VSS.n2173 272.089
R1844 VSS.n3418 VSS.n3392 272.089
R1845 VSS.n3415 VSS.n3414 272.089
R1846 VSS.n3418 VSS.n3391 272.089
R1847 VSS.n3415 VSS.n3396 272.089
R1848 VSS.n3418 VSS.n3390 272.089
R1849 VSS.n3415 VSS.n3395 272.089
R1850 VSS.n3418 VSS.n3389 272.089
R1851 VSS.n3415 VSS.n3394 272.089
R1852 VSS.n3418 VSS.n3388 272.089
R1853 VSS.n3416 VSS.n3415 272.089
R1854 VSS.n3933 VSS.n3922 272.089
R1855 VSS.n3931 VSS.n3923 272.089
R1856 VSS.n3935 VSS.n3923 272.089
R1857 VSS.n3928 VSS.n3922 272.089
R1858 VSS.n3940 VSS.n3923 272.089
R1859 VSS.n3942 VSS.n3922 272.089
R1860 VSS.n3944 VSS.n3923 272.089
R1861 VSS.n3925 VSS.n3922 272.089
R1862 VSS.n3949 VSS.n3923 272.089
R1863 VSS.n3951 VSS.n3922 272.089
R1864 VSS.n3953 VSS.n3923 272.089
R1865 VSS.n5074 VSS.n5073 272.089
R1866 VSS.n5084 VSS.n5055 272.089
R1867 VSS.n5074 VSS.n5062 272.089
R1868 VSS.n5084 VSS.n5056 272.089
R1869 VSS.n5074 VSS.n5061 272.089
R1870 VSS.n5084 VSS.n5057 272.089
R1871 VSS.n5076 VSS.n5074 272.089
R1872 VSS.n5084 VSS.n5058 272.089
R1873 VSS.n5074 VSS.n5059 272.089
R1874 VSS.n5084 VSS.n5083 272.089
R1875 VSS.n4551 VSS.n4535 272.089
R1876 VSS.n4559 VSS.n4558 272.089
R1877 VSS.n4552 VSS.n4551 272.089
R1878 VSS.n4559 VSS.n4533 272.089
R1879 VSS.n4551 VSS.n4538 272.089
R1880 VSS.n4559 VSS.n4532 272.089
R1881 VSS.n4551 VSS.n4539 272.089
R1882 VSS.n4559 VSS.n4531 272.089
R1883 VSS.n4551 VSS.n4550 272.089
R1884 VSS.n4559 VSS.n4530 272.089
R1885 VSS.n4551 VSS.n4528 272.089
R1886 VSS.n2988 VSS.n2987 272.089
R1887 VSS.n2998 VSS.n2967 272.089
R1888 VSS.n2988 VSS.n2974 272.089
R1889 VSS.n2998 VSS.n2968 272.089
R1890 VSS.n2988 VSS.n2973 272.089
R1891 VSS.n2998 VSS.n2969 272.089
R1892 VSS.n2990 VSS.n2988 272.089
R1893 VSS.n2998 VSS.n2970 272.089
R1894 VSS.n2988 VSS.n2971 272.089
R1895 VSS.n2998 VSS.n2997 272.089
R1896 VSS.n2938 VSS.n2930 272.089
R1897 VSS.n2939 VSS.n2931 272.089
R1898 VSS.n2944 VSS.n2931 272.089
R1899 VSS.n2946 VSS.n2930 272.089
R1900 VSS.n2948 VSS.n2931 272.089
R1901 VSS.n2935 VSS.n2930 272.089
R1902 VSS.n2953 VSS.n2931 272.089
R1903 VSS.n2955 VSS.n2930 272.089
R1904 VSS.n2957 VSS.n2931 272.089
R1905 VSS.n2932 VSS.n2930 272.089
R1906 VSS.n2962 VSS.n2931 272.089
R1907 VSS.n2118 VSS.n1841 272.089
R1908 VSS.n2119 VSS.n1841 272.089
R1909 VSS.n2133 VSS.n1841 272.089
R1910 VSS.n2134 VSS.n1841 272.089
R1911 VSS.n3971 VSS.n1841 272.089
R1912 VSS.n2146 VSS.n1841 272.089
R1913 VSS.n3203 VSS.n1841 272.089
R1914 VSS.n3341 VSS.n1841 272.089
R1915 VSS.n3209 VSS.n1841 272.089
R1916 VSS.n3225 VSS.n1841 272.089
R1917 VSS.n3226 VSS.n1841 272.089
R1918 VSS.n3311 VSS.n1841 272.089
R1919 VSS.n3920 VSS.n1841 272.089
R1920 VSS.n2219 VSS.n1841 272.089
R1921 VSS.n2345 VSS.n1841 272.089
R1922 VSS.n2344 VSS.n1841 272.089
R1923 VSS.n2331 VSS.n1841 272.089
R1924 VSS.n3442 VSS.n1841 272.089
R1925 VSS.n2328 VSS.n1841 272.089
R1926 VSS.n4594 VSS.n1841 272.089
R1927 VSS.n1845 VSS.n1841 272.089
R1928 VSS.n1861 VSS.n1841 272.089
R1929 VSS.n1862 VSS.n1841 272.089
R1930 VSS.n4564 VSS.n1841 272.089
R1931 VSS.n1915 VSS.n1841 272.089
R1932 VSS.n1888 VSS.n1844 272.089
R1933 VSS.n4575 VSS.n1844 272.089
R1934 VSS.n1858 VSS.n1844 272.089
R1935 VSS.n4592 VSS.n1844 272.089
R1936 VSS.n1844 VSS.n1840 272.089
R1937 VSS.n3440 VSS.n1844 272.089
R1938 VSS.n2373 VSS.n1844 272.089
R1939 VSS.n2364 VSS.n1844 272.089
R1940 VSS.n2355 VSS.n1844 272.089
R1941 VSS.n3918 VSS.n1844 272.089
R1942 VSS.n3310 VSS.n1844 272.089
R1943 VSS.n3322 VSS.n1844 272.089
R1944 VSS.n3222 VSS.n1844 272.089
R1945 VSS.n3339 VSS.n1844 272.089
R1946 VSS.n3206 VSS.n1844 272.089
R1947 VSS.n3969 VSS.n1844 272.089
R1948 VSS.n2143 VSS.n1844 272.089
R1949 VSS.n3982 VSS.n1844 272.089
R1950 VSS.n2131 VSS.n1844 272.089
R1951 VSS.n3995 VSS.n1844 272.089
R1952 VSS.n2758 VSS.n1748 272.089
R1953 VSS.n2754 VSS.n1743 272.089
R1954 VSS.n2763 VSS.n1748 272.089
R1955 VSS.n2765 VSS.n1743 272.089
R1956 VSS.n2767 VSS.n1748 272.089
R1957 VSS.n2751 VSS.n1743 272.089
R1958 VSS.n2772 VSS.n1748 272.089
R1959 VSS.n2774 VSS.n1743 272.089
R1960 VSS.n2750 VSS.n1748 272.089
R1961 VSS.n3004 VSS.n1744 272.089
R1962 VSS.n2816 VSS.n1752 272.089
R1963 VSS.n3009 VSS.n1744 272.089
R1964 VSS.n3011 VSS.n1752 272.089
R1965 VSS.n3013 VSS.n1744 272.089
R1966 VSS.n2813 VSS.n1752 272.089
R1967 VSS.n3018 VSS.n1744 272.089
R1968 VSS.n3020 VSS.n1752 272.089
R1969 VSS.n2812 VSS.n1744 272.089
R1970 VSS.n1991 VSS.n1745 272.089
R1971 VSS.n4515 VSS.n1749 272.089
R1972 VSS.n4513 VSS.n1745 272.089
R1973 VSS.n1993 VSS.n1749 272.089
R1974 VSS.n4508 VSS.n1745 272.089
R1975 VSS.n4506 VSS.n1749 272.089
R1976 VSS.n1995 VSS.n1745 272.089
R1977 VSS.n4501 VSS.n1749 272.089
R1978 VSS.n4499 VSS.n1745 272.089
R1979 VSS.n1984 VSS.n1953 272.089
R1980 VSS.n4525 VSS.n1957 272.089
R1981 VSS.n1984 VSS.n1983 272.089
R1982 VSS.n4525 VSS.n1958 272.089
R1983 VSS.n1984 VSS.n1968 272.089
R1984 VSS.n4525 VSS.n1959 272.089
R1985 VSS.n1984 VSS.n1967 272.089
R1986 VSS.n4525 VSS.n1960 272.089
R1987 VSS.n1986 VSS.n1984 272.089
R1988 VSS.n4525 VSS.n1961 272.089
R1989 VSS.n2695 VSS.n2694 272.089
R1990 VSS.n2778 VSS.n1743 272.089
R1991 VSS.n3024 VSS.n1752 272.089
R1992 VSS.n1997 VSS.n1749 272.089
R1993 VSS.n2756 VSS.n1743 272.089
R1994 VSS.n3002 VSS.n1752 272.089
R1995 VSS.n4520 VSS.n1749 272.089
R1996 VSS.n4687 VSS.n1700 272.089
R1997 VSS.n4687 VSS.n1699 272.089
R1998 VSS.n4687 VSS.n1698 272.089
R1999 VSS.n4687 VSS.n1697 272.089
R2000 VSS.n4687 VSS.n1696 272.089
R2001 VSS.n4687 VSS.n1694 272.089
R2002 VSS.n4687 VSS.n1693 272.089
R2003 VSS.n4687 VSS.n1692 272.089
R2004 VSS.n4687 VSS.n1691 272.089
R2005 VSS.n4687 VSS.n1690 272.089
R2006 VSS.n4687 VSS.n1688 272.089
R2007 VSS.n4687 VSS.n1687 272.089
R2008 VSS.n4687 VSS.n1686 272.089
R2009 VSS.n4687 VSS.n1685 272.089
R2010 VSS.n4687 VSS.n1684 272.089
R2011 VSS.n4687 VSS.n1682 272.089
R2012 VSS.n4687 VSS.n1681 272.089
R2013 VSS.n4687 VSS.n1680 272.089
R2014 VSS.n4687 VSS.n1679 272.089
R2015 VSS.n4687 VSS.n1678 272.089
R2016 VSS.n4688 VSS.n4687 272.089
R2017 VSS.n4687 VSS.n1676 272.089
R2018 VSS.n4687 VSS.n1675 272.089
R2019 VSS.n4687 VSS.n1674 272.089
R2020 VSS.n4687 VSS.n1673 272.089
R2021 VSS.n1826 VSS.n1707 272.089
R2022 VSS.n1826 VSS.n1825 272.089
R2023 VSS.n1826 VSS.n1785 272.089
R2024 VSS.n1826 VSS.n1784 272.089
R2025 VSS.n1826 VSS.n1783 272.089
R2026 VSS.n1826 VSS.n1670 272.089
R2027 VSS.n4430 VSS.n1826 272.089
R2028 VSS.n4423 VSS.n1826 272.089
R2029 VSS.n4414 VSS.n1826 272.089
R2030 VSS.n4405 VSS.n1826 272.089
R2031 VSS.n4624 VSS.n1826 272.089
R2032 VSS.n2923 VSS.n1826 272.089
R2033 VSS.n2898 VSS.n1826 272.089
R2034 VSS.n2891 VSS.n1826 272.089
R2035 VSS.n2882 VSS.n1826 272.089
R2036 VSS.n2873 VSS.n1826 272.089
R2037 VSS.n2864 VSS.n1826 272.089
R2038 VSS.n2393 VSS.n1826 272.089
R2039 VSS.n3380 VSS.n1826 272.089
R2040 VSS.n3264 VSS.n1826 272.089
R2041 VSS.n3255 VSS.n1826 272.089
R2042 VSS.n3246 VSS.n1826 272.089
R2043 VSS.n3371 VSS.n1826 272.089
R2044 VSS.n3190 VSS.n1826 272.089
R2045 VSS.n3148 VSS.n1826 272.089
R2046 VSS.n2559 VSS.n1826 272.089
R2047 VSS.n2549 VSS.n1826 272.089
R2048 VSS.n2572 VSS.n1826 272.089
R2049 VSS.n2537 VSS.n1826 272.089
R2050 VSS.n4007 VSS.n1826 272.089
R2051 VSS.n3155 VSS.n3154 272.089
R2052 VSS.n3415 VSS.n3387 272.089
R2053 VSS.n2988 VSS.n2929 272.089
R2054 VSS.n1984 VSS.n1963 272.089
R2055 VSS.n1949 VSS.n1841 272.089
R2056 VSS.n1945 VSS.n1841 272.089
R2057 VSS.n1893 VSS.n1841 272.089
R2058 VSS.n1931 VSS.n1841 272.089
R2059 VSS.n1906 VSS.n1841 272.089
R2060 VSS.n1917 VSS.n1844 272.089
R2061 VSS.n1929 VSS.n1844 272.089
R2062 VSS.n1904 VSS.n1844 272.089
R2063 VSS.n1943 VSS.n1844 272.089
R2064 VSS.n1947 VSS.n1844 272.089
R2065 VSS.n5410 VSS.n129 272.089
R2066 VSS.n131 VSS.n129 272.089
R2067 VSS.n139 VSS.n129 272.089
R2068 VSS.n140 VSS.n129 272.089
R2069 VSS.n155 VSS.n129 272.089
R2070 VSS.n5117 VSS.n129 272.089
R2071 VSS.n631 VSS.n129 272.089
R2072 VSS.n639 VSS.n129 272.089
R2073 VSS.n640 VSS.n129 272.089
R2074 VSS.n655 VSS.n129 272.089
R2075 VSS.n2245 VSS.n129 272.089
R2076 VSS.n2246 VSS.n129 272.089
R2077 VSS.n3471 VSS.n129 272.089
R2078 VSS.n3487 VSS.n129 272.089
R2079 VSS.n3507 VSS.n129 272.089
R2080 VSS.n4889 VSS.n129 272.089
R2081 VSS.n838 VSS.n129 272.089
R2082 VSS.n846 VSS.n129 272.089
R2083 VSS.n847 VSS.n129 272.089
R2084 VSS.n862 VSS.n129 272.089
R2085 VSS.n1278 VSS.n129 272.089
R2086 VSS.n1279 VSS.n129 272.089
R2087 VSS.n1424 VSS.n129 272.089
R2088 VSS.n1428 VSS.n129 272.089
R2089 VSS.n1409 VSS.n129 272.089
R2090 VSS.n1483 VSS.n130 272.089
R2091 VSS.n1426 VSS.n130 272.089
R2092 VSS.n1430 VSS.n130 272.089
R2093 VSS.n1415 VSS.n130 272.089
R2094 VSS.n4769 VSS.n130 272.089
R2095 VSS.n4740 VSS.n130 272.089
R2096 VSS.n4861 VSS.n130 272.089
R2097 VSS.n860 VSS.n130 272.089
R2098 VSS.n4874 VSS.n130 272.089
R2099 VSS.n844 VSS.n130 272.089
R2100 VSS.n4887 VSS.n130 272.089
R2101 VSS.n4891 VSS.n130 272.089
R2102 VSS.n3508 VSS.n130 272.089
R2103 VSS.n3466 VSS.n130 272.089
R2104 VSS.n3485 VSS.n130 272.089
R2105 VSS.n3476 VSS.n130 272.089
R2106 VSS.n3907 VSS.n130 272.089
R2107 VSS.n2420 VSS.n130 272.089
R2108 VSS.n5089 VSS.n130 272.089
R2109 VSS.n653 VSS.n130 272.089
R2110 VSS.n5102 VSS.n130 272.089
R2111 VSS.n637 VSS.n130 272.089
R2112 VSS.n5115 VSS.n130 272.089
R2113 VSS.n5119 VSS.n130 272.089
R2114 VSS.n5382 VSS.n130 272.089
R2115 VSS.n153 VSS.n130 272.089
R2116 VSS.n5395 VSS.n130 272.089
R2117 VSS.n137 VSS.n130 272.089
R2118 VSS.n5408 VSS.n130 272.089
R2119 VSS.n5412 VSS.n130 272.089
R2120 VSS.n5367 VSS.n161 272.089
R2121 VSS.n5074 VSS.n661 272.089
R2122 VSS.n5037 VSS.n674 272.089
R2123 VSS.n4846 VSS.n867 272.089
R2124 VSS.n1008 VSS.n272 272.089
R2125 VSS.n5003 VSS.n5002 272.089
R2126 VSS.n3645 VSS.n3644 272.089
R2127 VSS.n492 VSS.n243 272.089
R2128 VSS.n4228 VSS.n4227 270.175
R2129 VSS.n4784 VSS.n1233 264.301
R2130 VSS.n4784 VSS.n1244 264.301
R2131 VSS.n4108 VSS.n13 264.301
R2132 VSS.n4012 VSS.n2080 264.301
R2133 VSS.n4224 VSS.n127 264.301
R2134 VSS.n4198 VSS.n4073 264.301
R2135 VSS.n4134 VSS.n4133 264.301
R2136 VSS.n4684 VSS.n1728 264.301
R2137 VSS.n1487 VSS.n1486 264.301
R2138 VSS.n4333 VSS.n2054 259.416
R2139 VSS.n4721 VSS.n4720 258.334
R2140 VSS.n2020 VSS.n2019 258.334
R2141 VSS.n4631 VSS.n1760 258.334
R2142 VSS.n2794 VSS.n2793 258.334
R2143 VSS.n3090 VSS.n3089 258.334
R2144 VSS.n2439 VSS.n2224 258.334
R2145 VSS.n3433 VSS.n2391 258.334
R2146 VSS.n5436 VSS.n99 258.334
R2147 VSS.n5479 VSS.n5477 258.334
R2148 VSS.n5456 VSS.n60 258.334
R2149 VSS.n5178 VSS.n335 258.334
R2150 VSS.n5161 VSS.n364 258.334
R2151 VSS.n5143 VSS.n395 258.334
R2152 VSS.n1185 VSS.n1184 258.334
R2153 VSS.n4834 VSS.n892 258.334
R2154 VSS.n4762 VSS.n4761 258.334
R2155 VSS.n4958 VSS.n4956 258.334
R2156 VSS.n4933 VSS.n746 258.334
R2157 VSS.n4915 VSS.n780 258.334
R2158 VSS.n3830 VSS.n3829 258.334
R2159 VSS.n3865 VSS.n3864 258.334
R2160 VSS.n3900 VSS.n3899 258.334
R2161 VSS.n2116 VSS.n123 258.334
R2162 VSS.n4005 VSS.n2084 258.334
R2163 VSS.n3200 VSS.n419 258.334
R2164 VSS.n3364 VSS.n3363 258.334
R2165 VSS.n1837 VSS.n804 258.334
R2166 VSS.n4617 VSS.n4616 258.334
R2167 VSS.n3126 VSS.n3125 258.334
R2168 VSS.n5500 VSS.n6 254.34
R2169 VSS.n5502 VSS.n6 254.34
R2170 VSS.n5512 VSS.n6 254.34
R2171 VSS.n484 VSS.n6 254.34
R2172 VSS.n490 VSS.n6 254.34
R2173 VSS.n495 VSS.n6 254.34
R2174 VSS.n328 VSS.n6 254.34
R2175 VSS.n5202 VSS.n6 254.34
R2176 VSS.n5204 VSS.n6 254.34
R2177 VSS.n5217 VSS.n6 254.34
R2178 VSS.n5219 VSS.n6 254.34
R2179 VSS.n5233 VSS.n6 254.34
R2180 VSS.n5236 VSS.n6 254.34
R2181 VSS.n5248 VSS.n6 254.34
R2182 VSS.n5250 VSS.n6 254.34
R2183 VSS.n5263 VSS.n6 254.34
R2184 VSS.n5265 VSS.n6 254.34
R2185 VSS.n5279 VSS.n6 254.34
R2186 VSS.n5282 VSS.n6 254.34
R2187 VSS.n5294 VSS.n6 254.34
R2188 VSS.n5296 VSS.n6 254.34
R2189 VSS.n5309 VSS.n6 254.34
R2190 VSS.n5311 VSS.n6 254.34
R2191 VSS.n5325 VSS.n6 254.34
R2192 VSS.n1206 VSS.n6 254.34
R2193 VSS.n4816 VSS.n6 254.34
R2194 VSS.n1210 VSS.n6 254.34
R2195 VSS.n4804 VSS.n6 254.34
R2196 VSS.n1216 VSS.n6 254.34
R2197 VSS.n4791 VSS.n6 254.34
R2198 VSS.n2623 VSS.n2622 254.34
R2199 VSS.n4012 VSS.n2079 254.34
R2200 VSS.n4063 VSS.n127 254.34
R2201 VSS.n4078 VSS.n4073 254.34
R2202 VSS.n4133 VSS.n4131 254.34
R2203 VSS.n4332 VSS.n4321 254.34
R2204 VSS.n4684 VSS.n1727 254.34
R2205 VSS.n4784 VSS.n1226 254.34
R2206 VSS.n4784 VSS.n1225 254.34
R2207 VSS.n4784 VSS.n1224 254.34
R2208 VSS.n4784 VSS.n1223 254.34
R2209 VSS.n4784 VSS.n1222 254.34
R2210 VSS.n4784 VSS.n1232 254.34
R2211 VSS.n4784 VSS.n1231 254.34
R2212 VSS.n4784 VSS.n1230 254.34
R2213 VSS.n4784 VSS.n1229 254.34
R2214 VSS.n1487 VSS.n1408 254.34
R2215 VSS.n4784 VSS.n1228 254.34
R2216 VSS.n4784 VSS.n1246 254.34
R2217 VSS.n4784 VSS.n1238 254.34
R2218 VSS.n4784 VSS.n1237 254.34
R2219 VSS.n4784 VSS.n1236 254.34
R2220 VSS.n4784 VSS.n1235 254.34
R2221 VSS.n4784 VSS.n1234 254.34
R2222 VSS.n4785 VSS.n4784 254.34
R2223 VSS.n4784 VSS.n1243 254.34
R2224 VSS.n4784 VSS.n1242 254.34
R2225 VSS.n4784 VSS.n1241 254.34
R2226 VSS.n4784 VSS.n1240 254.34
R2227 VSS.n4302 VSS.n4301 252.179
R2228 VSS.n1724 VSS.n1627 250
R2229 VSS.n2051 VSS.n1650 250
R2230 VSS.n4451 VSS.n1765 250
R2231 VSS.n2818 VSS.n2403 250
R2232 VSS.n2744 VSS.n2472 250
R2233 VSS.n3447 VSS.n2228 250
R2234 VSS.n2852 VSS.n2851 250
R2235 VSS.n439 VSS.n438 250
R2236 VSS.n516 VSS.n515 250
R2237 VSS.n559 VSS.n558 250
R2238 VSS.n3729 VSS.n3728 250
R2239 VSS.n3732 VSS.n3731 250
R2240 VSS.n1339 VSS.n922 250
R2241 VSS.n1101 VSS.n1085 250
R2242 VSS.n1104 VSS.n1103 250
R2243 VSS.n3609 VSS.n2296 250
R2244 VSS.n3513 VSS.n2321 250
R2245 VSS.n2167 VSS.n109 250
R2246 VSS.n2517 VSS.n2516 250
R2247 VSS.n3306 VSS.n405 250
R2248 VSS.n3272 VSS.n3271 250
R2249 VSS.n1884 VSS.n790 250
R2250 VSS.n4393 VSS.n4392 250
R2251 VSS.n2657 VSS.n2524 250
R2252 VSS.n2625 VSS.n2589 249.663
R2253 VSS.n4110 VSS.t32 244.445
R2254 VSS.n4266 VSS.n4265 243.201
R2255 VSS.n4281 VSS.n4280 243.201
R2256 VSS.n4313 VSS.n4312 237.494
R2257 VSS.n4282 VSS.n4252 236.8
R2258 VSS.n4262 VSS.n4251 236.8
R2259 VSS.n4297 VSS.n4296 234
R2260 VSS.n4233 VSS.t79 229.225
R2261 VSS.n4233 VSS.t67 228.215
R2262 VSS.n4234 VSS.t83 228.215
R2263 VSS.n4235 VSS.t78 228.215
R2264 VSS.n4302 VSS.t88 225.507
R2265 VSS.n4717 VSS.n1623 221.667
R2266 VSS.n4228 VSS.t32 212.281
R2267 VSS.t35 VSS.n2628 207.214
R2268 VSS.t35 VSS.n2715 207.214
R2269 VSS.t35 VSS.n2802 207.214
R2270 VSS.n4468 VSS.t35 207.214
R2271 VSS.t35 VSS.n2028 207.214
R2272 VSS.n4275 VSS.n4268 201.927
R2273 VSS.n4790 VSS.n1218 197
R2274 VSS.n3110 VSS.t35 189.579
R2275 VSS.n3075 VSS.t35 189.579
R2276 VSS.n3040 VSS.t35 189.579
R2277 VSS.t35 VSS.n4456 189.579
R2278 VSS.n4348 VSS.t35 189.579
R2279 VSS.n5499 VSS.n12 187.249
R2280 VSS.t35 VSS.n1741 186.55
R2281 VSS.n4025 VSS.t32 186.55
R2282 VSS.n4053 VSS.t32 186.55
R2283 VSS.n4210 VSS.t32 186.55
R2284 VSS.n4146 VSS.t32 186.55
R2285 VSS.n4119 VSS.t32 186.55
R2286 VSS.n4310 VSS.n4231 185.225
R2287 VSS.n1709 VSS.n1253 185
R2288 VSS.n1711 VSS.n1710 185
R2289 VSS.n1713 VSS.n1712 185
R2290 VSS.n1715 VSS.n1714 185
R2291 VSS.n1717 VSS.n1716 185
R2292 VSS.n1719 VSS.n1718 185
R2293 VSS.n1721 VSS.n1720 185
R2294 VSS.n1723 VSS.n1722 185
R2295 VSS.n1725 VSS.n1724 185
R2296 VSS.n2036 VSS.n2035 185
R2297 VSS.n2038 VSS.n2037 185
R2298 VSS.n2040 VSS.n2039 185
R2299 VSS.n2042 VSS.n2041 185
R2300 VSS.n2044 VSS.n2043 185
R2301 VSS.n2046 VSS.n2045 185
R2302 VSS.n2048 VSS.n2047 185
R2303 VSS.n2050 VSS.n2049 185
R2304 VSS.n2052 VSS.n2051 185
R2305 VSS.n2019 VSS.n2018 185
R2306 VSS.n2017 VSS.n2016 185
R2307 VSS.n2015 VSS.n2014 185
R2308 VSS.n2013 VSS.n2012 185
R2309 VSS.n2011 VSS.n2010 185
R2310 VSS.n2009 VSS.n2008 185
R2311 VSS.n2007 VSS.n2006 185
R2312 VSS.n1666 VSS.n1665 185
R2313 VSS.n4710 VSS.n4709 185
R2314 VSS.n4436 VSS.n4435 185
R2315 VSS.n4438 VSS.n4437 185
R2316 VSS.n4440 VSS.n4439 185
R2317 VSS.n4442 VSS.n4441 185
R2318 VSS.n4444 VSS.n4443 185
R2319 VSS.n4446 VSS.n4445 185
R2320 VSS.n4448 VSS.n4447 185
R2321 VSS.n4450 VSS.n4449 185
R2322 VSS.n4452 VSS.n4451 185
R2323 VSS.n1760 VSS.n1758 185
R2324 VSS.n2909 VSS.n2908 185
R2325 VSS.n2911 VSS.n2910 185
R2326 VSS.n2913 VSS.n2912 185
R2327 VSS.n2915 VSS.n2914 185
R2328 VSS.n2917 VSS.n2916 185
R2329 VSS.n2919 VSS.n2918 185
R2330 VSS.n2921 VSS.n2920 185
R2331 VSS.n2922 VSS.n1779 185
R2332 VSS.n2835 VSS.n2834 185
R2333 VSS.n2833 VSS.n2832 185
R2334 VSS.n2831 VSS.n2830 185
R2335 VSS.n2829 VSS.n2828 185
R2336 VSS.n2827 VSS.n2826 185
R2337 VSS.n2825 VSS.n2824 185
R2338 VSS.n2823 VSS.n2822 185
R2339 VSS.n2821 VSS.n2820 185
R2340 VSS.n2819 VSS.n2818 185
R2341 VSS.n2793 VSS.n2792 185
R2342 VSS.n2791 VSS.n2790 185
R2343 VSS.n2789 VSS.n2788 185
R2344 VSS.n2787 VSS.n2786 185
R2345 VSS.n2785 VSS.n2784 185
R2346 VSS.n2419 VSS.n2418 185
R2347 VSS.n3427 VSS.n3426 185
R2348 VSS.n3425 VSS.n2417 185
R2349 VSS.n3424 VSS.n3423 185
R2350 VSS.n2468 VSS.n2464 185
R2351 VSS.n2731 VSS.n2730 185
R2352 VSS.n2733 VSS.n2732 185
R2353 VSS.n2735 VSS.n2734 185
R2354 VSS.n2737 VSS.n2736 185
R2355 VSS.n2739 VSS.n2738 185
R2356 VSS.n2741 VSS.n2740 185
R2357 VSS.n2743 VSS.n2742 185
R2358 VSS.n2745 VSS.n2744 185
R2359 VSS.n3089 VSS.n2712 185
R2360 VSS.n2711 VSS.n2710 185
R2361 VSS.n2709 VSS.n2708 185
R2362 VSS.n2707 VSS.n2706 185
R2363 VSS.n2705 VSS.n2704 185
R2364 VSS.n2703 VSS.n2702 185
R2365 VSS.n2701 VSS.n2700 185
R2366 VSS.n2699 VSS.n2698 185
R2367 VSS.n2493 VSS.n2486 185
R2368 VSS.n2440 VSS.n2439 185
R2369 VSS.n2438 VSS.n2437 185
R2370 VSS.n2436 VSS.n2435 185
R2371 VSS.n2434 VSS.n2433 185
R2372 VSS.n2432 VSS.n2431 185
R2373 VSS.n2430 VSS.n2429 185
R2374 VSS.n2428 VSS.n2427 185
R2375 VSS.n2426 VSS.n2425 185
R2376 VSS.n2424 VSS.n2242 185
R2377 VSS.n2458 VSS.n2391 185
R2378 VSS.n2457 VSS.n2456 185
R2379 VSS.n2455 VSS.n2454 185
R2380 VSS.n2453 VSS.n2452 185
R2381 VSS.n2451 VSS.n2450 185
R2382 VSS.n2449 VSS.n2448 185
R2383 VSS.n2447 VSS.n2446 185
R2384 VSS.n2445 VSS.n2444 185
R2385 VSS.n2443 VSS.n2442 185
R2386 VSS.n2334 VSS.n2322 185
R2387 VSS.n2837 VSS.n2836 185
R2388 VSS.n2839 VSS.n2838 185
R2389 VSS.n2841 VSS.n2840 185
R2390 VSS.n2843 VSS.n2842 185
R2391 VSS.n2845 VSS.n2844 185
R2392 VSS.n2847 VSS.n2846 185
R2393 VSS.n2849 VSS.n2848 185
R2394 VSS.n2851 VSS.n2850 185
R2395 VSS.n3464 VSS.n3463 185
R2396 VSS.n3462 VSS.n3461 185
R2397 VSS.n3460 VSS.n3459 185
R2398 VSS.n3458 VSS.n3457 185
R2399 VSS.n3456 VSS.n3455 185
R2400 VSS.n3454 VSS.n3453 185
R2401 VSS.n3452 VSS.n3451 185
R2402 VSS.n3450 VSS.n3449 185
R2403 VSS.n3448 VSS.n3447 185
R2404 VSS.n126 VSS.n99 185
R2405 VSS.n4175 VSS.n4174 185
R2406 VSS.n4177 VSS.n4176 185
R2407 VSS.n4179 VSS.n4178 185
R2408 VSS.n4181 VSS.n4180 185
R2409 VSS.n4183 VSS.n4182 185
R2410 VSS.n4185 VSS.n4184 185
R2411 VSS.n4187 VSS.n4186 185
R2412 VSS.n4189 VSS.n4188 185
R2413 VSS.n456 VSS.n455 185
R2414 VSS.n454 VSS.n453 185
R2415 VSS.n452 VSS.n451 185
R2416 VSS.n450 VSS.n449 185
R2417 VSS.n448 VSS.n447 185
R2418 VSS.n446 VSS.n445 185
R2419 VSS.n444 VSS.n443 185
R2420 VSS.n442 VSS.n441 185
R2421 VSS.n440 VSS.n439 185
R2422 VSS.n5480 VSS.n5479 185
R2423 VSS.n5481 VSS.n17 185
R2424 VSS.n5483 VSS.n5482 185
R2425 VSS.n5485 VSS.n16 185
R2426 VSS.n5488 VSS.n5487 185
R2427 VSS.n5489 VSS.n15 185
R2428 VSS.n5491 VSS.n5490 185
R2429 VSS.n5493 VSS.n14 185
R2430 VSS.n5496 VSS.n5495 185
R2431 VSS.n4173 VSS.n60 185
R2432 VSS.n4172 VSS.n4171 185
R2433 VSS.n4170 VSS.n4169 185
R2434 VSS.n4168 VSS.n4167 185
R2435 VSS.n4166 VSS.n4165 185
R2436 VSS.n4164 VSS.n4163 185
R2437 VSS.n4162 VSS.n4161 185
R2438 VSS.n4160 VSS.n4159 185
R2439 VSS.n4158 VSS.n4157 185
R2440 VSS.n526 VSS.n525 185
R2441 VSS.n528 VSS.n527 185
R2442 VSS.n530 VSS.n529 185
R2443 VSS.n532 VSS.n531 185
R2444 VSS.n534 VSS.n533 185
R2445 VSS.n536 VSS.n535 185
R2446 VSS.n538 VSS.n537 185
R2447 VSS.n540 VSS.n539 185
R2448 VSS.n558 VSS.n541 185
R2449 VSS.n501 VSS.n478 185
R2450 VSS.n503 VSS.n502 185
R2451 VSS.n504 VSS.n477 185
R2452 VSS.n506 VSS.n505 185
R2453 VSS.n508 VSS.n475 185
R2454 VSS.n510 VSS.n509 185
R2455 VSS.n511 VSS.n474 185
R2456 VSS.n513 VSS.n512 185
R2457 VSS.n515 VSS.n457 185
R2458 VSS.n517 VSS.n516 185
R2459 VSS.n516 VSS.t40 185
R2460 VSS.n473 VSS.n471 185
R2461 VSS.n462 VSS.n38 185
R2462 VSS.n5461 VSS.n5460 185
R2463 VSS.n5464 VSS.n5463 185
R2464 VSS.n37 VSS.n33 185
R2465 VSS.n35 VSS.n25 185
R2466 VSS.n34 VSS.n24 185
R2467 VSS.n5477 VSS.n5476 185
R2468 VSS.n459 VSS.n458 185
R2469 VSS.n461 VSS.n50 185
R2470 VSS.t62 VSS.n50 185
R2471 VSS.n463 VSS.n41 185
R2472 VSS.n5459 VSS.n5458 185
R2473 VSS.n40 VSS.n32 185
R2474 VSS.n46 VSS.n31 185
R2475 VSS.n45 VSS.n44 185
R2476 VSS.n5473 VSS.n5472 185
R2477 VSS.n5475 VSS.n5474 185
R2478 VSS.n560 VSS.n559 185
R2479 VSS.n556 VSS.n555 185
R2480 VSS.n554 VSS.n553 185
R2481 VSS.n5441 VSS.n5440 185
R2482 VSS.n5443 VSS.n5442 185
R2483 VSS.n75 VSS.n74 185
R2484 VSS.n73 VSS.n67 185
R2485 VSS.n66 VSS.n61 185
R2486 VSS.n5456 VSS.n5455 185
R2487 VSS.t62 VSS.n5456 185
R2488 VSS.n543 VSS.n542 185
R2489 VSS.n557 VSS.n89 185
R2490 VSS.t36 VSS.n89 185
R2491 VSS.n552 VSS.n80 185
R2492 VSS.n5439 VSS.n5438 185
R2493 VSS.n79 VSS.n77 185
R2494 VSS.n85 VSS.n76 185
R2495 VSS.n84 VSS.n83 185
R2496 VSS.n5452 VSS.n5451 185
R2497 VSS.n5454 VSS.n5453 185
R2498 VSS.n5229 VSS.n5228 185
R2499 VSS.n317 VSS.n316 185
R2500 VSS.n3717 VSS.n3716 185
R2501 VSS.n3719 VSS.n3718 185
R2502 VSS.n3721 VSS.n3713 185
R2503 VSS.n3723 VSS.n3722 185
R2504 VSS.n3724 VSS.n3712 185
R2505 VSS.n3726 VSS.n3725 185
R2506 VSS.n3728 VSS.n3711 185
R2507 VSS.n437 VSS.n364 185
R2508 VSS.n436 VSS.n435 185
R2509 VSS.n434 VSS.n433 185
R2510 VSS.n432 VSS.n431 185
R2511 VSS.n430 VSS.n429 185
R2512 VSS.n428 VSS.n427 185
R2513 VSS.n426 VSS.n425 185
R2514 VSS.n424 VSS.n423 185
R2515 VSS.n422 VSS.n336 185
R2516 VSS.n5178 VSS.n5177 185
R2517 VSS.n5180 VSS.n334 185
R2518 VSS.n5183 VSS.n5182 185
R2519 VSS.n5184 VSS.n333 185
R2520 VSS.n5186 VSS.n5185 185
R2521 VSS.n5188 VSS.n332 185
R2522 VSS.n5191 VSS.n5190 185
R2523 VSS.n5192 VSS.n331 185
R2524 VSS.n5195 VSS.n5194 185
R2525 VSS.n3730 VSS.n3729 185
R2526 VSS.n3729 VSS.t50 185
R2527 VSS.n3710 VSS.n3673 185
R2528 VSS.n3708 VSS.n3707 185
R2529 VSS.n3693 VSS.n3674 185
R2530 VSS.n3688 VSS.n3687 185
R2531 VSS.n3685 VSS.n3684 185
R2532 VSS.n5167 VSS.n5166 185
R2533 VSS.n5170 VSS.n5169 185
R2534 VSS.n337 VSS.n335 185
R2535 VSS.n3801 VSS.n3800 185
R2536 VSS.n3704 VSS.n3703 185
R2537 VSS.n3706 VSS.n3705 185
R2538 VSS.n3692 VSS.n3691 185
R2539 VSS.n3690 VSS.n3689 185
R2540 VSS.n3683 VSS.n344 185
R2541 VSS.n5165 VSS.n5164 185
R2542 VSS.n345 VSS.n340 185
R2543 VSS.n357 VSS.n339 185
R2544 VSS.n629 VSS.n395 185
R2545 VSS.n628 VSS.n627 185
R2546 VSS.n626 VSS.n625 185
R2547 VSS.n624 VSS.n623 185
R2548 VSS.n622 VSS.n621 185
R2549 VSS.n620 VSS.n619 185
R2550 VSS.n618 VSS.n617 185
R2551 VSS.n616 VSS.n615 185
R2552 VSS.n614 VSS.n613 185
R2553 VSS.n3749 VSS.n3748 185
R2554 VSS.n3747 VSS.n3746 185
R2555 VSS.n3745 VSS.n3744 185
R2556 VSS.n3743 VSS.n3742 185
R2557 VSS.n3741 VSS.n3740 185
R2558 VSS.n3739 VSS.n3738 185
R2559 VSS.n3737 VSS.n3736 185
R2560 VSS.n3735 VSS.n3734 185
R2561 VSS.n3733 VSS.n3732 185
R2562 VSS.n3799 VSS.n3798 185
R2563 VSS.n3797 VSS.n3796 185
R2564 VSS.n3795 VSS.n3794 185
R2565 VSS.n3793 VSS.n3792 185
R2566 VSS.n3791 VSS.n3790 185
R2567 VSS.n3789 VSS.n3788 185
R2568 VSS.n3787 VSS.n3786 185
R2569 VSS.n3785 VSS.n3784 185
R2570 VSS.n3783 VSS.n3782 185
R2571 VSS.n1186 VSS.n1185 185
R2572 VSS.n1188 VSS.n1187 185
R2573 VSS.n1190 VSS.n1189 185
R2574 VSS.n1192 VSS.n1191 185
R2575 VSS.n1194 VSS.n1193 185
R2576 VSS.n1196 VSS.n1195 185
R2577 VSS.n1198 VSS.n1197 185
R2578 VSS.n1200 VSS.n1199 185
R2579 VSS.n1201 VSS.n937 185
R2580 VSS.n4761 VSS.n4760 185
R2581 VSS.n4759 VSS.n4758 185
R2582 VSS.n4757 VSS.n4756 185
R2583 VSS.n4755 VSS.n4754 185
R2584 VSS.n4753 VSS.n4752 185
R2585 VSS.n4751 VSS.n4750 185
R2586 VSS.n4749 VSS.n4748 185
R2587 VSS.n4747 VSS.n4746 185
R2588 VSS.n4745 VSS.n4744 185
R2589 VSS.n938 VSS.n892 185
R2590 VSS.n940 VSS.n939 185
R2591 VSS.n942 VSS.n941 185
R2592 VSS.n944 VSS.n943 185
R2593 VSS.n946 VSS.n945 185
R2594 VSS.n948 VSS.n947 185
R2595 VSS.n950 VSS.n949 185
R2596 VSS.n952 VSS.n951 185
R2597 VSS.n953 VSS.n910 185
R2598 VSS.n1589 VSS.n1588 185
R2599 VSS.n1587 VSS.n1586 185
R2600 VSS.n1310 VSS.n1309 185
R2601 VSS.n1308 VSS.n1307 185
R2602 VSS.n1604 VSS.n1603 185
R2603 VSS.n1602 VSS.n1601 185
R2604 VSS.n1297 VSS.n1296 185
R2605 VSS.n1295 VSS.n893 185
R2606 VSS.n4835 VSS.n4834 185
R2607 VSS.n1585 VSS.n1584 185
R2608 VSS.n1319 VSS.n1318 185
R2609 VSS.n1317 VSS.n1316 185
R2610 VSS.n1598 VSS.n1597 185
R2611 VSS.n1600 VSS.n1599 185
R2612 VSS.n1306 VSS.n1305 185
R2613 VSS.n1304 VSS.n1303 185
R2614 VSS.n1613 VSS.n1612 185
R2615 VSS.n1614 VSS.n891 185
R2616 VSS.n1564 VSS.n1563 185
R2617 VSS.n1566 VSS.n1565 185
R2618 VSS.n1568 VSS.n1567 185
R2619 VSS.n1570 VSS.n1569 185
R2620 VSS.n1572 VSS.n1571 185
R2621 VSS.n1574 VSS.n1573 185
R2622 VSS.n1576 VSS.n1575 185
R2623 VSS.n1578 VSS.n1577 185
R2624 VSS.n1580 VSS.n1579 185
R2625 VSS.n1324 VSS.n1323 185
R2626 VSS.n1326 VSS.n1325 185
R2627 VSS.n1328 VSS.n1327 185
R2628 VSS.n1330 VSS.n1329 185
R2629 VSS.n1332 VSS.n1331 185
R2630 VSS.n1334 VSS.n1333 185
R2631 VSS.n1336 VSS.n1335 185
R2632 VSS.n1338 VSS.n1337 185
R2633 VSS.n1340 VSS.n1339 185
R2634 VSS.n1342 VSS.n922 185
R2635 VSS.t53 VSS.n922 185
R2636 VSS.n1345 VSS.n1344 185
R2637 VSS.n1348 VSS.n1346 185
R2638 VSS.n1350 VSS.n1349 185
R2639 VSS.n1352 VSS.n1351 185
R2640 VSS.n1356 VSS.n919 185
R2641 VSS.n4824 VSS.n4823 185
R2642 VSS.n918 VSS.n913 185
R2643 VSS.n1184 VSS.n912 185
R2644 VSS.n1562 VSS.n1561 185
R2645 VSS.n1377 VSS.n1376 185
R2646 VSS.n1375 VSS.n1374 185
R2647 VSS.n1368 VSS.n1367 185
R2648 VSS.n1366 VSS.n1365 185
R2649 VSS.n1359 VSS.n1358 185
R2650 VSS.n1357 VSS.n917 185
R2651 VSS.n916 VSS.n911 185
R2652 VSS.n4831 VSS.n4830 185
R2653 VSS.n5321 VSS.n5320 185
R2654 VSS.n279 VSS.n278 185
R2655 VSS.n1091 VSS.n1088 185
R2656 VSS.n1093 VSS.n1092 185
R2657 VSS.n1094 VSS.n1087 185
R2658 VSS.n1096 VSS.n1095 185
R2659 VSS.n1098 VSS.n1086 185
R2660 VSS.n1099 VSS.n1037 185
R2661 VSS.n1102 VSS.n1101 185
R2662 VSS.n819 VSS.n746 185
R2663 VSS.n818 VSS.n817 185
R2664 VSS.n816 VSS.n815 185
R2665 VSS.n814 VSS.n813 185
R2666 VSS.n812 VSS.n811 185
R2667 VSS.n810 VSS.n809 185
R2668 VSS.n808 VSS.n807 185
R2669 VSS.n726 VSS.n725 185
R2670 VSS.n4937 VSS.n4936 185
R2671 VSS.n4956 VSS.n4939 185
R2672 VSS.n4954 VSS.n4953 185
R2673 VSS.n4952 VSS.n4940 185
R2674 VSS.n4951 VSS.n4950 185
R2675 VSS.n4948 VSS.n4941 185
R2676 VSS.n4946 VSS.n4945 185
R2677 VSS.n4944 VSS.n4943 185
R2678 VSS.n292 VSS.n291 185
R2679 VSS.n5287 VSS.n5286 185
R2680 VSS.n1085 VSS.n1084 185
R2681 VSS.n1085 VSS.t51 185
R2682 VSS.n1078 VSS.n1038 185
R2683 VSS.n1074 VSS.n1073 185
R2684 VSS.n1071 VSS.n1042 185
R2685 VSS.n1069 VSS.n1068 185
R2686 VSS.n1054 VSS.n1044 185
R2687 VSS.n1049 VSS.n724 185
R2688 VSS.n4961 VSS.n4960 185
R2689 VSS.n4958 VSS.n4957 185
R2690 VSS.n1170 VSS.n1036 185
R2691 VSS.n1075 VSS.n1039 185
R2692 VSS.n1077 VSS.n1076 185
R2693 VSS.n1065 VSS.n1064 185
R2694 VSS.n1067 VSS.n1066 185
R2695 VSS.n1053 VSS.n1052 185
R2696 VSS.n1051 VSS.n1050 185
R2697 VSS.n728 VSS.n723 185
R2698 VSS.n727 VSS.n722 185
R2699 VSS.n837 VSS.n780 185
R2700 VSS.n836 VSS.n835 185
R2701 VSS.n834 VSS.n833 185
R2702 VSS.n832 VSS.n831 185
R2703 VSS.n830 VSS.n829 185
R2704 VSS.n828 VSS.n827 185
R2705 VSS.n826 VSS.n825 185
R2706 VSS.n824 VSS.n823 185
R2707 VSS.n822 VSS.n821 185
R2708 VSS.n1121 VSS.n1120 185
R2709 VSS.n1119 VSS.n1118 185
R2710 VSS.n1117 VSS.n1116 185
R2711 VSS.n1115 VSS.n1114 185
R2712 VSS.n1113 VSS.n1112 185
R2713 VSS.n1111 VSS.n1110 185
R2714 VSS.n1109 VSS.n1108 185
R2715 VSS.n1107 VSS.n1106 185
R2716 VSS.n1105 VSS.n1104 185
R2717 VSS.n1172 VSS.n1171 185
R2718 VSS.n1169 VSS.n1168 185
R2719 VSS.n1167 VSS.n1166 185
R2720 VSS.n1165 VSS.n1164 185
R2721 VSS.n1163 VSS.n1162 185
R2722 VSS.n1161 VSS.n1160 185
R2723 VSS.n1159 VSS.n1158 185
R2724 VSS.n1157 VSS.n1156 185
R2725 VSS.n1155 VSS.n1154 185
R2726 VSS.n1146 VSS.n1145 185
R2727 VSS.n1144 VSS.n1143 185
R2728 VSS.n1137 VSS.n1136 185
R2729 VSS.n1135 VSS.n1134 185
R2730 VSS.n4920 VSS.n4919 185
R2731 VSS.n4922 VSS.n4921 185
R2732 VSS.n753 VSS.n752 185
R2733 VSS.n751 VSS.n745 185
R2734 VSS.n4933 VSS.n4932 185
R2735 VSS.n1123 VSS.n1122 185
R2736 VSS.n1125 VSS.n770 185
R2737 VSS.t46 VSS.n770 185
R2738 VSS.n1127 VSS.n1126 185
R2739 VSS.n1129 VSS.n762 185
R2740 VSS.n4918 VSS.n4917 185
R2741 VSS.n764 VSS.n760 185
R2742 VSS.n763 VSS.n759 185
R2743 VSS.n4929 VSS.n4928 185
R2744 VSS.n4931 VSS.n4930 185
R2745 VSS.n5275 VSS.n5274 185
R2746 VSS.n298 VSS.n297 185
R2747 VSS.n3589 VSS.n3586 185
R2748 VSS.n3591 VSS.n3590 185
R2749 VSS.n3592 VSS.n3585 185
R2750 VSS.n3594 VSS.n3593 185
R2751 VSS.n3596 VSS.n3583 185
R2752 VSS.n3598 VSS.n3597 185
R2753 VSS.n3599 VSS.n2296 185
R2754 VSS.n3864 VSS.n2269 185
R2755 VSS.n3862 VSS.n3861 185
R2756 VSS.n3860 VSS.n2270 185
R2757 VSS.n3859 VSS.n3858 185
R2758 VSS.n3856 VSS.n2271 185
R2759 VSS.n3854 VSS.n3853 185
R2760 VSS.n3852 VSS.n2272 185
R2761 VSS.n3851 VSS.n3850 185
R2762 VSS.n3848 VSS.n2273 185
R2763 VSS.n3829 VSS.n3812 185
R2764 VSS.n3827 VSS.n3826 185
R2765 VSS.n3825 VSS.n3813 185
R2766 VSS.n3824 VSS.n3823 185
R2767 VSS.n3821 VSS.n3814 185
R2768 VSS.n3819 VSS.n3818 185
R2769 VSS.n3817 VSS.n3816 185
R2770 VSS.n311 VSS.n310 185
R2771 VSS.n5241 VSS.n5240 185
R2772 VSS.n3609 VSS.n3608 185
R2773 VSS.n3609 VSS.t57 185
R2774 VSS.n3614 VSS.n3613 185
R2775 VSS.n3611 VSS.n2287 185
R2776 VSS.n3610 VSS.n2286 185
R2777 VSS.n3629 VSS.n3628 185
R2778 VSS.n3837 VSS.n3836 185
R2779 VSS.n3834 VSS.n3833 185
R2780 VSS.n3832 VSS.n2276 185
R2781 VSS.n3830 VSS.n2275 185
R2782 VSS.n3607 VSS.n3606 185
R2783 VSS.n3604 VSS.n2295 185
R2784 VSS.n3603 VSS.n2294 185
R2785 VSS.n3621 VSS.n3620 185
R2786 VSS.n3627 VSS.n3626 185
R2787 VSS.n3624 VSS.n2282 185
R2788 VSS.n3623 VSS.n2281 185
R2789 VSS.n2278 VSS.n2274 185
R2790 VSS.n3846 VSS.n3845 185
R2791 VSS.n3899 VSS.n2251 185
R2792 VSS.n3897 VSS.n3896 185
R2793 VSS.n3895 VSS.n2252 185
R2794 VSS.n3894 VSS.n3893 185
R2795 VSS.n3891 VSS.n2253 185
R2796 VSS.n3889 VSS.n3888 185
R2797 VSS.n3887 VSS.n2254 185
R2798 VSS.n3886 VSS.n3885 185
R2799 VSS.n3883 VSS.n2255 185
R2800 VSS.n3528 VSS.n2308 185
R2801 VSS.n3527 VSS.n3526 185
R2802 VSS.n3525 VSS.n3524 185
R2803 VSS.n3523 VSS.n2318 185
R2804 VSS.n3521 VSS.n3520 185
R2805 VSS.n3519 VSS.n2319 185
R2806 VSS.n3518 VSS.n3517 185
R2807 VSS.n3515 VSS.n2320 185
R2808 VSS.n3513 VSS.n3512 185
R2809 VSS.n3602 VSS.n3601 185
R2810 VSS.n3582 VSS.n3581 185
R2811 VSS.n3580 VSS.n2304 185
R2812 VSS.n3578 VSS.n3577 185
R2813 VSS.n3576 VSS.n2305 185
R2814 VSS.n3575 VSS.n3574 185
R2815 VSS.n3572 VSS.n2306 185
R2816 VSS.n3570 VSS.n3569 185
R2817 VSS.n3568 VSS.n2307 185
R2818 VSS.n3560 VSS.n3559 185
R2819 VSS.n3557 VSS.n2312 185
R2820 VSS.n3555 VSS.n3554 185
R2821 VSS.n3548 VSS.n2314 185
R2822 VSS.n3538 VSS.n2265 185
R2823 VSS.n3872 VSS.n3871 185
R2824 VSS.n3869 VSS.n3868 185
R2825 VSS.n3867 VSS.n2258 185
R2826 VSS.n3865 VSS.n2257 185
R2827 VSS.n3530 VSS.n2309 185
R2828 VSS.n3531 VSS.n2311 185
R2829 VSS.n3531 VSS.t59 185
R2830 VSS.n3553 VSS.n3552 185
R2831 VSS.n3550 VSS.n3549 185
R2832 VSS.n3537 VSS.n3536 185
R2833 VSS.n3534 VSS.n2264 185
R2834 VSS.n3533 VSS.n2263 185
R2835 VSS.n2260 VSS.n2256 185
R2836 VSS.n3881 VSS.n3880 185
R2837 VSS.n3774 VSS.n3773 185
R2838 VSS.n3772 VSS.n3771 185
R2839 VSS.n3765 VSS.n3764 185
R2840 VSS.n3763 VSS.n3762 185
R2841 VSS.n5148 VSS.n5147 185
R2842 VSS.n5150 VSS.n5149 185
R2843 VSS.n371 VSS.n370 185
R2844 VSS.n369 VSS.n363 185
R2845 VSS.n5161 VSS.n5160 185
R2846 VSS.n3751 VSS.n3750 185
R2847 VSS.n3753 VSS.n385 185
R2848 VSS.t63 VSS.n385 185
R2849 VSS.n3755 VSS.n3754 185
R2850 VSS.n3757 VSS.n377 185
R2851 VSS.n5146 VSS.n5145 185
R2852 VSS.n379 VSS.n375 185
R2853 VSS.n378 VSS.n374 185
R2854 VSS.n5157 VSS.n5156 185
R2855 VSS.n5159 VSS.n5158 185
R2856 VSS.n125 VSS.n123 185
R2857 VSS.n5430 VSS.n5429 185
R2858 VSS.n5428 VSS.n124 185
R2859 VSS.n5427 VSS.n5426 185
R2860 VSS.n5425 VSS.n5424 185
R2861 VSS.n5423 VSS.n5422 185
R2862 VSS.n5421 VSS.n5420 185
R2863 VSS.n5419 VSS.n5418 185
R2864 VSS.n5417 VSS.n5416 185
R2865 VSS.n2084 VSS.n2081 185
R2866 VSS.n2106 VSS.n2105 185
R2867 VSS.n2108 VSS.n2107 185
R2868 VSS.n2110 VSS.n2109 185
R2869 VSS.n2112 VSS.n2111 185
R2870 VSS.n2113 VSS.n2104 185
R2871 VSS.n4003 VSS.n4002 185
R2872 VSS.n4001 VSS.n2103 185
R2873 VSS.n4000 VSS.n3999 185
R2874 VSS.n2499 VSS.n2150 185
R2875 VSS.n2501 VSS.n2500 185
R2876 VSS.n2503 VSS.n2502 185
R2877 VSS.n2505 VSS.n2504 185
R2878 VSS.n2507 VSS.n2506 185
R2879 VSS.n2509 VSS.n2508 185
R2880 VSS.n2511 VSS.n2510 185
R2881 VSS.n2513 VSS.n2512 185
R2882 VSS.n2516 VSS.n2514 185
R2883 VSS.n2152 VSS.n2151 185
R2884 VSS.n2154 VSS.n2153 185
R2885 VSS.n2156 VSS.n2155 185
R2886 VSS.n2158 VSS.n2157 185
R2887 VSS.n2160 VSS.n2159 185
R2888 VSS.n2162 VSS.n2161 185
R2889 VSS.n2164 VSS.n2163 185
R2890 VSS.n2166 VSS.n2165 185
R2891 VSS.n2168 VSS.n2167 185
R2892 VSS.n421 VSS.n419 185
R2893 VSS.n5137 VSS.n5136 185
R2894 VSS.n5135 VSS.n420 185
R2895 VSS.n5134 VSS.n5133 185
R2896 VSS.n5132 VSS.n5131 185
R2897 VSS.n5130 VSS.n5129 185
R2898 VSS.n5128 VSS.n5127 185
R2899 VSS.n5126 VSS.n5125 185
R2900 VSS.n5124 VSS.n5123 185
R2901 VSS.n3363 VSS.n3194 185
R2902 VSS.n3361 VSS.n3360 185
R2903 VSS.n3359 VSS.n3195 185
R2904 VSS.n3358 VSS.n3357 185
R2905 VSS.n3355 VSS.n3196 185
R2906 VSS.n3353 VSS.n3352 185
R2907 VSS.n3351 VSS.n3197 185
R2908 VSS.n3350 VSS.n3349 185
R2909 VSS.n3347 VSS.n3198 185
R2910 VSS.n3289 VSS.n3288 185
R2911 VSS.n3287 VSS.n3232 185
R2912 VSS.n3285 VSS.n3284 185
R2913 VSS.n3283 VSS.n3233 185
R2914 VSS.n3282 VSS.n3281 185
R2915 VSS.n3279 VSS.n3234 185
R2916 VSS.n3277 VSS.n3276 185
R2917 VSS.n3275 VSS.n3274 185
R2918 VSS.n3272 VSS.n2465 185
R2919 VSS.n3291 VSS.n3290 185
R2920 VSS.n3293 VSS.n3292 185
R2921 VSS.n3295 VSS.n3294 185
R2922 VSS.n3297 VSS.n3296 185
R2923 VSS.n3299 VSS.n3298 185
R2924 VSS.n3301 VSS.n3300 185
R2925 VSS.n3303 VSS.n3302 185
R2926 VSS.n3305 VSS.n3304 185
R2927 VSS.n3307 VSS.n3306 185
R2928 VSS.n3231 VSS.n405 185
R2929 VSS.t56 VSS.n405 185
R2930 VSS.n3319 VSS.n3318 185
R2931 VSS.n3220 VSS.n3219 185
R2932 VSS.n3218 VSS.n3217 185
R2933 VSS.n3334 VSS.n3333 185
R2934 VSS.n3336 VSS.n3335 185
R2935 VSS.n3212 VSS.n3211 185
R2936 VSS.n3210 VSS.n3202 185
R2937 VSS.n3201 VSS.n3200 185
R2938 VSS.n3315 VSS.n3314 185
R2939 VSS.n3317 VSS.n3316 185
R2940 VSS.n3316 VSS.t49 185
R2941 VSS.n3229 VSS.n3227 185
R2942 VSS.n3326 VSS.n3325 185
R2943 VSS.n3332 VSS.n3331 185
R2944 VSS.n3329 VSS.n3214 185
R2945 VSS.n3328 VSS.n3213 185
R2946 VSS.n3207 VSS.n3199 185
R2947 VSS.n3345 VSS.n3344 185
R2948 VSS.n2147 VSS.n109 185
R2949 VSS.t31 VSS.n109 185
R2950 VSS.n2141 VSS.n2140 185
R2951 VSS.n3977 VSS.n3976 185
R2952 VSS.n3979 VSS.n3978 185
R2953 VSS.n2129 VSS.n2128 185
R2954 VSS.n2127 VSS.n2126 185
R2955 VSS.n3990 VSS.n3989 185
R2956 VSS.n3992 VSS.n3991 185
R2957 VSS.n2117 VSS.n2116 185
R2958 VSS.n2149 VSS.n2148 185
R2959 VSS.n2144 VSS.n2093 185
R2960 VSS.t54 VSS.n2093 185
R2961 VSS.n3975 VSS.n3974 185
R2962 VSS.n2138 VSS.n2137 185
R2963 VSS.n2136 VSS.n2135 185
R2964 VSS.n3986 VSS.n3985 185
R2965 VSS.n3988 VSS.n3987 185
R2966 VSS.n2123 VSS.n2122 185
R2967 VSS.n2121 VSS.n2120 185
R2968 VSS.n806 VSS.n804 185
R2969 VSS.n4909 VSS.n4908 185
R2970 VSS.n4907 VSS.n805 185
R2971 VSS.n4906 VSS.n4905 185
R2972 VSS.n4904 VSS.n4903 185
R2973 VSS.n4902 VSS.n4901 185
R2974 VSS.n4900 VSS.n4899 185
R2975 VSS.n4898 VSS.n4897 185
R2976 VSS.n4896 VSS.n4895 185
R2977 VSS.n4616 VSS.n1831 185
R2978 VSS.n4614 VSS.n4613 185
R2979 VSS.n4612 VSS.n1832 185
R2980 VSS.n4611 VSS.n4610 185
R2981 VSS.n4608 VSS.n1833 185
R2982 VSS.n4606 VSS.n4605 185
R2983 VSS.n4604 VSS.n1834 185
R2984 VSS.n4603 VSS.n4602 185
R2985 VSS.n4600 VSS.n1835 185
R2986 VSS.n4378 VSS.n4376 185
R2987 VSS.n4380 VSS.n4379 185
R2988 VSS.n4381 VSS.n4375 185
R2989 VSS.n4383 VSS.n4382 185
R2990 VSS.n4385 VSS.n4373 185
R2991 VSS.n4387 VSS.n4386 185
R2992 VSS.n4388 VSS.n4372 185
R2993 VSS.n4390 VSS.n4389 185
R2994 VSS.n4392 VSS.n4367 185
R2995 VSS.n1869 VSS.n1868 185
R2996 VSS.n1871 VSS.n1870 185
R2997 VSS.n1873 VSS.n1872 185
R2998 VSS.n1875 VSS.n1874 185
R2999 VSS.n1877 VSS.n1876 185
R3000 VSS.n1879 VSS.n1878 185
R3001 VSS.n1881 VSS.n1880 185
R3002 VSS.n1883 VSS.n1882 185
R3003 VSS.n1885 VSS.n1884 185
R3004 VSS.n1867 VSS.n790 185
R3005 VSS.t43 VSS.n790 185
R3006 VSS.n4572 VSS.n4571 185
R3007 VSS.n1856 VSS.n1855 185
R3008 VSS.n1854 VSS.n1853 185
R3009 VSS.n4587 VSS.n4586 185
R3010 VSS.n4589 VSS.n4588 185
R3011 VSS.n1848 VSS.n1847 185
R3012 VSS.n1846 VSS.n1839 185
R3013 VSS.n1838 VSS.n1837 185
R3014 VSS.n4568 VSS.n4567 185
R3015 VSS.n4570 VSS.n4569 185
R3016 VSS.n4569 VSS.t33 185
R3017 VSS.n1865 VSS.n1863 185
R3018 VSS.n4579 VSS.n4578 185
R3019 VSS.n4585 VSS.n4584 185
R3020 VSS.n4582 VSS.n1850 185
R3021 VSS.n4581 VSS.n1849 185
R3022 VSS.n1842 VSS.n1836 185
R3023 VSS.n4598 VSS.n4597 185
R3024 VSS.n3437 VSS.n2228 185
R3025 VSS.t65 VSS.n2228 185
R3026 VSS.n2343 VSS.n2342 185
R3027 VSS.n2367 VSS.n2341 185
R3028 VSS.n2369 VSS.n2368 185
R3029 VSS.n2361 VSS.n2360 185
R3030 VSS.n2359 VSS.n2358 185
R3031 VSS.n2352 VSS.n2222 185
R3032 VSS.n3915 VSS.n3914 185
R3033 VSS.n2224 VSS.n2223 185
R3034 VSS.n3436 VSS.n3435 185
R3035 VSS.n2333 VSS.n2332 185
R3036 VSS.t47 VSS.n2333 185
R3037 VSS.n2377 VSS.n2376 185
R3038 VSS.n2370 VSS.n2340 185
R3039 VSS.n2348 VSS.n2347 185
R3040 VSS.n2349 VSS.n2346 185
R3041 VSS.n2351 VSS.n2350 185
R3042 VSS.n2384 VSS.n2221 185
R3043 VSS.n2385 VSS.n2220 185
R3044 VSS.n2520 VSS.n2515 185
R3045 VSS.n2644 VSS.n2643 185
R3046 VSS.n2646 VSS.n2645 185
R3047 VSS.n2648 VSS.n2647 185
R3048 VSS.n2650 VSS.n2649 185
R3049 VSS.n2652 VSS.n2651 185
R3050 VSS.n2654 VSS.n2653 185
R3051 VSS.n2656 VSS.n2655 185
R3052 VSS.n2658 VSS.n2657 185
R3053 VSS.n3127 VSS.n3126 185
R3054 VSS.n3129 VSS.n3128 185
R3055 VSS.n3131 VSS.n3130 185
R3056 VSS.n3133 VSS.n3132 185
R3057 VSS.n3135 VSS.n3134 185
R3058 VSS.n3137 VSS.n3136 185
R3059 VSS.n3139 VSS.n3138 185
R3060 VSS.n3141 VSS.n3140 185
R3061 VSS.n3142 VSS.n2082 185
R3062 VSS.n3102 VSS.n2524 185
R3063 VSS.t34 VSS.n2524 185
R3064 VSS.n3105 VSS.n3104 185
R3065 VSS.n2642 VSS.n2641 185
R3066 VSS.n2640 VSS.n2635 185
R3067 VSS.n3114 VSS.n3113 185
R3068 VSS.n3116 VSS.n3115 185
R3069 VSS.n2633 VSS.n2632 185
R3070 VSS.n2631 VSS.n2585 185
R3071 VSS.n3125 VSS.n3124 185
R3072 VSS.n3067 VSS.n2472 185
R3073 VSS.t64 VSS.n2472 185
R3074 VSS.n3070 VSS.n3069 185
R3075 VSS.n2729 VSS.n2728 185
R3076 VSS.n2727 VSS.n2722 185
R3077 VSS.n3079 VSS.n3078 185
R3078 VSS.n3081 VSS.n3080 185
R3079 VSS.n2720 VSS.n2719 185
R3080 VSS.n2718 VSS.n2713 185
R3081 VSS.n3091 VSS.n3090 185
R3082 VSS.n3032 VSS.n2403 185
R3083 VSS.t61 VSS.n2403 185
R3084 VSS.n3035 VSS.n3034 185
R3085 VSS.n2808 VSS.n2807 185
R3086 VSS.n2806 VSS.n2799 185
R3087 VSS.n3044 VSS.n3043 185
R3088 VSS.n3046 VSS.n3045 185
R3089 VSS.n3050 VSS.n3049 185
R3090 VSS.n3048 VSS.n2797 185
R3091 VSS.n2795 VSS.n2794 185
R3092 VSS.n4490 VSS.n1765 185
R3093 VSS.t44 VSS.n1765 185
R3094 VSS.n4454 VSS.n4453 185
R3095 VSS.n4481 VSS.n4480 185
R3096 VSS.n4479 VSS.n4477 185
R3097 VSS.n4475 VSS.n4474 185
R3098 VSS.n4473 VSS.n4472 185
R3099 VSS.n4460 VSS.n4459 185
R3100 VSS.n4461 VSS.n1761 185
R3101 VSS.n4632 VSS.n4631 185
R3102 VSS.n4340 VSS.n1650 185
R3103 VSS.t58 VSS.n1650 185
R3104 VSS.n4343 VSS.n4342 185
R3105 VSS.n2034 VSS.n2033 185
R3106 VSS.n2032 VSS.n2025 185
R3107 VSS.n4352 VSS.n4351 185
R3108 VSS.n4354 VSS.n4353 185
R3109 VSS.n4358 VSS.n4357 185
R3110 VSS.n4356 VSS.n2023 185
R3111 VSS.n2021 VSS.n2020 185
R3112 VSS.n2518 VSS.n2517 185
R3113 VSS.n2555 VSS.n2554 185
R3114 VSS.n2553 VSS.n2552 185
R3115 VSS.n2567 VSS.n2566 185
R3116 VSS.n2569 VSS.n2568 185
R3117 VSS.n2543 VSS.n2542 185
R3118 VSS.n2541 VSS.n2540 185
R3119 VSS.n2534 VSS.n2085 185
R3120 VSS.n4006 VSS.n4005 185
R3121 VSS.n4005 VSS.t54 185
R3122 VSS.n3271 VSS.n2466 185
R3123 VSS.n3269 VSS.n3268 185
R3124 VSS.n3236 VSS.n3235 185
R3125 VSS.n3239 VSS.n3237 185
R3126 VSS.n3242 VSS.n3241 185
R3127 VSS.n3243 VSS.n2492 185
R3128 VSS.n3368 VSS.n3367 185
R3129 VSS.n3365 VSS.n2488 185
R3130 VSS.n3364 VSS.n2487 185
R3131 VSS.n3364 VSS.t49 185
R3132 VSS.n2853 VSS.n2852 185
R3133 VSS.n2855 VSS.n2854 185
R3134 VSS.n2857 VSS.n2856 185
R3135 VSS.n2859 VSS.n2858 185
R3136 VSS.n2861 VSS.n2860 185
R3137 VSS.n2867 VSS.n2862 185
R3138 VSS.n2869 VSS.n2868 185
R3139 VSS.n2399 VSS.n2392 185
R3140 VSS.n3433 VSS.n3432 185
R3141 VSS.t47 VSS.n3433 185
R3142 VSS.n4393 VSS.n4368 185
R3143 VSS.n4395 VSS.n4369 185
R3144 VSS.n4396 VSS.n4370 185
R3145 VSS.n4398 VSS.n4371 185
R3146 VSS.n4401 VSS.n4400 185
R3147 VSS.n4402 VSS.n1830 185
R3148 VSS.n4621 VSS.n4620 185
R3149 VSS.n4618 VSS.n1781 185
R3150 VSS.n4617 VSS.n1780 185
R3151 VSS.n4617 VSS.t33 185
R3152 VSS.n1822 VSS.n1627 185
R3153 VSS.t48 VSS.n1627 185
R3154 VSS.n1815 VSS.n1814 185
R3155 VSS.n1804 VSS.n1787 185
R3156 VSS.n1806 VSS.n1805 185
R3157 VSS.n1793 VSS.n1788 185
R3158 VSS.n1795 VSS.n1794 185
R3159 VSS.n1789 VSS.n1643 185
R3160 VSS.n4715 VSS.n4714 185
R3161 VSS.t48 VSS.n4715 185
R3162 VSS.n1669 VSS.n1642 185
R3163 VSS.n3147 VSS.n3146 185
R3164 VSS.n2556 VSS.n2519 185
R3165 VSS.n2563 VSS.n2562 185
R3166 VSS.n2565 VSS.n2564 185
R3167 VSS.n2546 VSS.n2545 185
R3168 VSS.n2544 VSS.n2532 185
R3169 VSS.n2576 VSS.n2575 185
R3170 VSS.n2533 VSS.n2521 185
R3171 VSS.t34 VSS.n2521 185
R3172 VSS.n3143 VSS.n2083 185
R3173 VSS.n3379 VSS.n3378 185
R3174 VSS.n3267 VSS.n2467 185
R3175 VSS.n3261 VSS.n3260 185
R3176 VSS.n3259 VSS.n3258 185
R3177 VSS.n3252 VSS.n3251 185
R3178 VSS.n3250 VSS.n3249 185
R3179 VSS.n2491 VSS.n2490 185
R3180 VSS.n2489 VSS.n2469 185
R3181 VSS.t64 VSS.n2469 185
R3182 VSS.n3375 VSS.n3374 185
R3183 VSS.n2897 VSS.n2896 185
R3184 VSS.n2895 VSS.n2894 185
R3185 VSS.n2888 VSS.n2887 185
R3186 VSS.n2886 VSS.n2885 185
R3187 VSS.n2879 VSS.n2878 185
R3188 VSS.n2877 VSS.n2876 185
R3189 VSS.n2870 VSS.n2398 185
R3190 VSS.n3429 VSS.n2400 185
R3191 VSS.n3429 VSS.t61 185
R3192 VSS.n3431 VSS.n3430 185
R3193 VSS.n4429 VSS.n4428 185
R3194 VSS.n4427 VSS.n4426 185
R3195 VSS.n4420 VSS.n4419 185
R3196 VSS.n4418 VSS.n4417 185
R3197 VSS.n4411 VSS.n4410 185
R3198 VSS.n4409 VSS.n4408 185
R3199 VSS.n1829 VSS.n1828 185
R3200 VSS.n1827 VSS.n1762 185
R3201 VSS.t44 VSS.n1762 185
R3202 VSS.n4628 VSS.n4627 185
R3203 VSS.n1821 VSS.n1820 185
R3204 VSS.n1819 VSS.n1816 185
R3205 VSS.n1812 VSS.n1811 185
R3206 VSS.n1810 VSS.n1809 185
R3207 VSS.n1801 VSS.n1800 185
R3208 VSS.n1799 VSS.n1798 185
R3209 VSS.n1790 VSS.n1647 185
R3210 VSS.n4713 VSS.n4712 185
R3211 VSS.n4712 VSS.t58 185
R3212 VSS.n1668 VSS.n1646 185
R3213 VSS.n4707 VSS.n4706 185
R3214 VSS.n4705 VSS.n4704 185
R3215 VSS.n4703 VSS.n4702 185
R3216 VSS.n4701 VSS.n4700 185
R3217 VSS.n4699 VSS.n4698 185
R3218 VSS.n4697 VSS.n4696 185
R3219 VSS.n4695 VSS.n4694 185
R3220 VSS.n4693 VSS.n4692 185
R3221 VSS.n4691 VSS.n1623 185
R3222 VSS.n4722 VSS.n4721 185
R3223 VSS.n4724 VSS.n4723 185
R3224 VSS.n4726 VSS.n4725 185
R3225 VSS.n4728 VSS.n4727 185
R3226 VSS.n4730 VSS.n4729 185
R3227 VSS.n4732 VSS.n4731 185
R3228 VSS.n4734 VSS.n4733 185
R3229 VSS.n4736 VSS.n4735 185
R3230 VSS.n4737 VSS.n1274 185
R3231 VSS.n1920 VSS.n1257 185
R3232 VSS.n1926 VSS.n1925 185
R3233 VSS.n1908 VSS.n1907 185
R3234 VSS.n1910 VSS.n1909 185
R3235 VSS.n1938 VSS.n1937 185
R3236 VSS.n1940 VSS.n1939 185
R3237 VSS.n1898 VSS.n1897 185
R3238 VSS.n1896 VSS.n1895 185
R3239 VSS.n4720 VSS.n4719 185
R3240 VSS.n1922 VSS.n1921 185
R3241 VSS.n1924 VSS.n1923 185
R3242 VSS.n1914 VSS.n1913 185
R3243 VSS.n1912 VSS.n1911 185
R3244 VSS.n1936 VSS.n1935 185
R3245 VSS.n1934 VSS.n1901 185
R3246 VSS.n1900 VSS.n1899 185
R3247 VSS.n1894 VSS.n1624 185
R3248 VSS.n4718 VSS.n4717 185
R3249 VSS.n1464 VSS.n1463 185
R3250 VSS.n1461 VSS.n1460 185
R3251 VSS.n1459 VSS.n1458 185
R3252 VSS.n1457 VSS.n1456 185
R3253 VSS.n1455 VSS.n1454 185
R3254 VSS.n1453 VSS.n1452 185
R3255 VSS.n1451 VSS.n1450 185
R3256 VSS.n1256 VSS.n1255 185
R3257 VSS.n4777 VSS.n4776 185
R3258 VSS.n1583 VSS.n1582 185
R3259 VSS.n1465 VSS.n1321 185
R3260 VSS.n1467 VSS.n1466 185
R3261 VSS.n1469 VSS.n1468 185
R3262 VSS.n1471 VSS.n1470 185
R3263 VSS.n1473 VSS.n1472 185
R3264 VSS.n1475 VSS.n1474 185
R3265 VSS.n1477 VSS.n1476 185
R3266 VSS.n1479 VSS.n1478 185
R3267 VSS.n438 VSS.n150 185
R3268 VSS.n5390 VSS.n5389 185
R3269 VSS.n5392 VSS.n5391 185
R3270 VSS.n143 VSS.n142 185
R3271 VSS.n141 VSS.n135 185
R3272 VSS.n5403 VSS.n5402 185
R3273 VSS.n5405 VSS.n5404 185
R3274 VSS.n105 VSS.n100 185
R3275 VSS.n5436 VSS.n5435 185
R3276 VSS.t36 VSS.n5436 185
R3277 VSS.n3731 VSS.n650 185
R3278 VSS.n5097 VSS.n5096 185
R3279 VSS.n5099 VSS.n5098 185
R3280 VSS.n643 VSS.n642 185
R3281 VSS.n641 VSS.n635 185
R3282 VSS.n5110 VSS.n5109 185
R3283 VSS.n5112 VSS.n5111 185
R3284 VSS.n401 VSS.n396 185
R3285 VSS.n5143 VSS.n5142 185
R3286 VSS.t63 VSS.n5143 185
R3287 VSS.n3504 VSS.n2321 185
R3288 VSS.n3500 VSS.n3499 185
R3289 VSS.n3497 VSS.n3468 185
R3290 VSS.n3495 VSS.n3494 185
R3291 VSS.n3472 VSS.n3470 185
R3292 VSS.n3473 VSS.n2250 185
R3293 VSS.n3904 VSS.n3903 185
R3294 VSS.n3901 VSS.n2244 185
R3295 VSS.n3900 VSS.n2243 185
R3296 VSS.n3900 VSS.t59 185
R3297 VSS.n1103 VSS.n857 185
R3298 VSS.n4869 VSS.n4868 185
R3299 VSS.n4871 VSS.n4870 185
R3300 VSS.n850 VSS.n849 185
R3301 VSS.n848 VSS.n842 185
R3302 VSS.n4882 VSS.n4881 185
R3303 VSS.n4884 VSS.n4883 185
R3304 VSS.n786 VSS.n781 185
R3305 VSS.n4915 VSS.n4914 185
R3306 VSS.t46 VSS.n4915 185
R3307 VSS.n1448 VSS.n1447 185
R3308 VSS.n1446 VSS.n1445 185
R3309 VSS.n1440 VSS.n1439 185
R3310 VSS.n1438 VSS.n1437 185
R3311 VSS.n1414 VSS.n1413 185
R3312 VSS.n1418 VSS.n1283 185
R3313 VSS.n4766 VSS.n4765 185
R3314 VSS.n1282 VSS.n1277 185
R3315 VSS.n4762 VSS.n1276 185
R3316 VSS.n5386 VSS.n5385 185
R3317 VSS.n5388 VSS.n5387 185
R3318 VSS.n147 VSS.n146 185
R3319 VSS.n145 VSS.n144 185
R3320 VSS.n5399 VSS.n5398 185
R3321 VSS.n5401 VSS.n5400 185
R3322 VSS.n132 VSS.n104 185
R3323 VSS.n5432 VSS.n106 185
R3324 VSS.n5432 VSS.t31 185
R3325 VSS.n5434 VSS.n5433 185
R3326 VSS.n5093 VSS.n5092 185
R3327 VSS.n5095 VSS.n5094 185
R3328 VSS.n647 VSS.n646 185
R3329 VSS.n645 VSS.n644 185
R3330 VSS.n5106 VSS.n5105 185
R3331 VSS.n5108 VSS.n5107 185
R3332 VSS.n632 VSS.n400 185
R3333 VSS.n5139 VSS.n402 185
R3334 VSS.n5139 VSS.t56 185
R3335 VSS.n5141 VSS.n5140 185
R3336 VSS.n3501 VSS.n3465 185
R3337 VSS.n3503 VSS.n3502 185
R3338 VSS.n3491 VSS.n3490 185
R3339 VSS.n3493 VSS.n3492 185
R3340 VSS.n3482 VSS.n3481 185
R3341 VSS.n3480 VSS.n3479 185
R3342 VSS.n2249 VSS.n2248 185
R3343 VSS.n2247 VSS.n2225 185
R3344 VSS.t65 VSS.n2225 185
R3345 VSS.n3911 VSS.n3910 185
R3346 VSS.n4865 VSS.n4864 185
R3347 VSS.n4867 VSS.n4866 185
R3348 VSS.n854 VSS.n853 185
R3349 VSS.n852 VSS.n851 185
R3350 VSS.n4878 VSS.n4877 185
R3351 VSS.n4880 VSS.n4879 185
R3352 VSS.n839 VSS.n785 185
R3353 VSS.n4911 VSS.n787 185
R3354 VSS.n4911 VSS.t43 185
R3355 VSS.n4913 VSS.n4912 185
R3356 VSS.n1462 VSS.n1449 185
R3357 VSS.n1444 VSS.n1443 185
R3358 VSS.n1442 VSS.n1441 185
R3359 VSS.n1436 VSS.n1435 185
R3360 VSS.n1434 VSS.n1433 185
R3361 VSS.n1421 VSS.n1420 185
R3362 VSS.n1419 VSS.n1281 185
R3363 VSS.n1280 VSS.n1275 185
R3364 VSS.n4773 VSS.n4772 185
R3365 VSS.n499 VSS.n498 185
R3366 VSS.n487 VSS.n481 185
R3367 VSS.n486 VSS.n2 185
R3368 VSS.n5519 VSS.n5518 185
R3369 VSS.n5516 VSS.n5515 185
R3370 VSS.n4 VSS.n3 185
R3371 VSS.n5509 VSS.n5508 185
R3372 VSS.n5506 VSS.n5505 185
R3373 VSS.n5506 VSS.t40 185
R3374 VSS.n10 VSS.n9 185
R3375 VSS.n5226 VSS.n315 185
R3376 VSS.n5225 VSS.n319 185
R3377 VSS.n5223 VSS.n5222 185
R3378 VSS.n5214 VSS.n320 185
R3379 VSS.n5213 VSS.n5212 185
R3380 VSS.n5210 VSS.n324 185
R3381 VSS.n5208 VSS.n5207 185
R3382 VSS.n5199 VSS.n325 185
R3383 VSS.n325 VSS.t50 185
R3384 VSS.n5198 VSS.n5197 185
R3385 VSS.n5272 VSS.n296 185
R3386 VSS.n5271 VSS.n300 185
R3387 VSS.n5269 VSS.n5268 185
R3388 VSS.n5260 VSS.n301 185
R3389 VSS.n5259 VSS.n5258 185
R3390 VSS.n5256 VSS.n305 185
R3391 VSS.n5254 VSS.n5253 185
R3392 VSS.n5245 VSS.n306 185
R3393 VSS.n306 VSS.t57 185
R3394 VSS.n5244 VSS.n5243 185
R3395 VSS.n5318 VSS.n277 185
R3396 VSS.n5317 VSS.n281 185
R3397 VSS.n5315 VSS.n5314 185
R3398 VSS.n5306 VSS.n282 185
R3399 VSS.n5305 VSS.n5304 185
R3400 VSS.n5302 VSS.n286 185
R3401 VSS.n5300 VSS.n5299 185
R3402 VSS.n5291 VSS.n287 185
R3403 VSS.n287 VSS.t51 185
R3404 VSS.n5290 VSS.n5289 185
R3405 VSS.n4795 VSS.n4794 185
R3406 VSS.n4797 VSS.n4796 185
R3407 VSS.n4801 VSS.n4800 185
R3408 VSS.n4799 VSS.n1213 185
R3409 VSS.n4808 VSS.n4807 185
R3410 VSS.n4810 VSS.n4809 185
R3411 VSS.n4813 VSS.n4812 185
R3412 VSS.n1205 VSS.n920 185
R3413 VSS.t53 VSS.n920 185
R3414 VSS.n4820 VSS.n4819 185
R3415 VSS.n1554 VSS.n1553 175.546
R3416 VSS.n1550 VSS.n1549 175.546
R3417 VSS.n1546 VSS.n1545 175.546
R3418 VSS.n1542 VSS.n1541 175.546
R3419 VSS.n1538 VSS.n1221 175.546
R3420 VSS.n4786 VSS.n1219 175.546
R3421 VSS.n1516 VSS.n1515 175.546
R3422 VSS.n1520 VSS.n1519 175.546
R3423 VSS.n1524 VSS.n1523 175.546
R3424 VSS.n1528 VSS.n1527 175.546
R3425 VSS.n1532 VSS.n1531 175.546
R3426 VSS.n1491 VSS.n1490 175.546
R3427 VSS.n1495 VSS.n1494 175.546
R3428 VSS.n1499 VSS.n1498 175.546
R3429 VSS.n1503 VSS.n1502 175.546
R3430 VSS.n1507 VSS.n1506 175.546
R3431 VSS.n1248 VSS.n1247 175.546
R3432 VSS.n1389 VSS.n1247 175.546
R3433 VSS.n1393 VSS.n1392 175.546
R3434 VSS.n1397 VSS.n1396 175.546
R3435 VSS.n1401 VSS.n1400 175.546
R3436 VSS.n1405 VSS.n1404 175.546
R3437 VSS.n4681 VSS.n4652 175.546
R3438 VSS.n4681 VSS.n4653 175.546
R3439 VSS.n4677 VSS.n4653 175.546
R3440 VSS.n4677 VSS.n4658 175.546
R3441 VSS.n4673 VSS.n4658 175.546
R3442 VSS.n4673 VSS.n4660 175.546
R3443 VSS.n4669 VSS.n4660 175.546
R3444 VSS.n4669 VSS.n4662 175.546
R3445 VSS.n4665 VSS.n4662 175.546
R3446 VSS.n4665 VSS.n1249 175.546
R3447 VSS.n4155 VSS.n4079 175.546
R3448 VSS.n4155 VSS.n4080 175.546
R3449 VSS.n4151 VSS.n4080 175.546
R3450 VSS.n4151 VSS.n4084 175.546
R3451 VSS.n4147 VSS.n4084 175.546
R3452 VSS.n4147 VSS.n4086 175.546
R3453 VSS.n4143 VSS.n4086 175.546
R3454 VSS.n4143 VSS.n4088 175.546
R3455 VSS.n4139 VSS.n4088 175.546
R3456 VSS.n4139 VSS.n4090 175.546
R3457 VSS.n4219 VSS.n4061 175.546
R3458 VSS.n4219 VSS.n4062 175.546
R3459 VSS.n4215 VSS.n4062 175.546
R3460 VSS.n4215 VSS.n4068 175.546
R3461 VSS.n4211 VSS.n4068 175.546
R3462 VSS.n4211 VSS.n4070 175.546
R3463 VSS.n4207 VSS.n4070 175.546
R3464 VSS.n4207 VSS.n4072 175.546
R3465 VSS.n4203 VSS.n4072 175.546
R3466 VSS.n4203 VSS.n4074 175.546
R3467 VSS.n4039 VSS.n2064 175.546
R3468 VSS.n4043 VSS.n2064 175.546
R3469 VSS.n4043 VSS.n2062 175.546
R3470 VSS.n4048 VSS.n2062 175.546
R3471 VSS.n4048 VSS.n2060 175.546
R3472 VSS.n4052 VSS.n2060 175.546
R3473 VSS.n4052 VSS.n2059 175.546
R3474 VSS.n4057 VSS.n2059 175.546
R3475 VSS.n4057 VSS.n2057 175.546
R3476 VSS.n4223 VSS.n2057 175.546
R3477 VSS.n4225 VSS.n4223 175.546
R3478 VSS.n4015 VSS.n2077 175.546
R3479 VSS.n4015 VSS.n2075 175.546
R3480 VSS.n4020 VSS.n2075 175.546
R3481 VSS.n4020 VSS.n2073 175.546
R3482 VSS.n4024 VSS.n2073 175.546
R3483 VSS.n4024 VSS.n2072 175.546
R3484 VSS.n4028 VSS.n2072 175.546
R3485 VSS.n4028 VSS.n2070 175.546
R3486 VSS.n4033 VSS.n2070 175.546
R3487 VSS.n4033 VSS.n2066 175.546
R3488 VSS.n4130 VSS.n4098 175.546
R3489 VSS.n4126 VSS.n4098 175.546
R3490 VSS.n4126 VSS.n4101 175.546
R3491 VSS.n4122 VSS.n4101 175.546
R3492 VSS.n4122 VSS.n4120 175.546
R3493 VSS.n4120 VSS.n4104 175.546
R3494 VSS.n4116 VSS.n4104 175.546
R3495 VSS.n4116 VSS.n4106 175.546
R3496 VSS.n4112 VSS.n4106 175.546
R3497 VSS.n4112 VSS.n4109 175.546
R3498 VSS.n2621 VSS.n2591 175.546
R3499 VSS.n2617 VSS.n2591 175.546
R3500 VSS.n2617 VSS.n2593 175.546
R3501 VSS.n2613 VSS.n2593 175.546
R3502 VSS.n2613 VSS.n2612 175.546
R3503 VSS.n2612 VSS.n2611 175.546
R3504 VSS.n2611 VSS.n2595 175.546
R3505 VSS.n2607 VSS.n2595 175.546
R3506 VSS.n2607 VSS.n2604 175.546
R3507 VSS.n2604 VSS.n2603 175.546
R3508 VSS.n2625 VSS.n2586 175.546
R3509 VSS.n3122 VSS.n2586 175.546
R3510 VSS.n3122 VSS.n2587 175.546
R3511 VSS.n3118 VSS.n2587 175.546
R3512 VSS.n3118 VSS.n2629 175.546
R3513 VSS.n3111 VSS.n2629 175.546
R3514 VSS.n3111 VSS.n2636 175.546
R3515 VSS.n3107 VSS.n2636 175.546
R3516 VSS.n3107 VSS.n2638 175.546
R3517 VSS.n3100 VSS.n2638 175.546
R3518 VSS.n3100 VSS.n2660 175.546
R3519 VSS.n5503 VSS.n5501 175.546
R3520 VSS.n5511 VSS.n7 175.546
R3521 VSS.n5513 VSS.n5 175.546
R3522 VSS.n489 VSS.n485 175.546
R3523 VSS.n496 VSS.n491 175.546
R3524 VSS.n4817 VSS.n1207 175.546
R3525 VSS.n4815 VSS.n1208 175.546
R3526 VSS.n4805 VSS.n1211 175.546
R3527 VSS.n4803 VSS.n1212 175.546
R3528 VSS.n4792 VSS.n1217 175.546
R3529 VSS.n5201 VSS.n329 175.546
R3530 VSS.n5205 VSS.n5203 175.546
R3531 VSS.n5216 VSS.n322 175.546
R3532 VSS.n5220 VSS.n5218 175.546
R3533 VSS.n5232 VSS.n314 175.546
R3534 VSS.n5293 VSS.n289 175.546
R3535 VSS.n5297 VSS.n5295 175.546
R3536 VSS.n5308 VSS.n284 175.546
R3537 VSS.n5312 VSS.n5310 175.546
R3538 VSS.n5324 VSS.n276 175.546
R3539 VSS.n5247 VSS.n308 175.546
R3540 VSS.n5251 VSS.n5249 175.546
R3541 VSS.n5262 VSS.n303 175.546
R3542 VSS.n5266 VSS.n5264 175.546
R3543 VSS.n5278 VSS.n295 175.546
R3544 VSS.n3095 VSS.n2664 175.546
R3545 VSS.n3087 VSS.n2664 175.546
R3546 VSS.n3087 VSS.n2714 175.546
R3547 VSS.n3083 VSS.n2714 175.546
R3548 VSS.n3083 VSS.n2716 175.546
R3549 VSS.n3076 VSS.n2716 175.546
R3550 VSS.n3076 VSS.n2723 175.546
R3551 VSS.n3072 VSS.n2723 175.546
R3552 VSS.n3072 VSS.n2725 175.546
R3553 VSS.n3065 VSS.n2725 175.546
R3554 VSS.n3065 VSS.n3063 175.546
R3555 VSS.n3057 VSS.n3056 175.546
R3556 VSS.n3056 VSS.n2780 175.546
R3557 VSS.n3052 VSS.n2780 175.546
R3558 VSS.n3052 VSS.n2783 175.546
R3559 VSS.n2800 VSS.n2783 175.546
R3560 VSS.n3041 VSS.n2800 175.546
R3561 VSS.n3041 VSS.n2801 175.546
R3562 VSS.n3037 VSS.n2801 175.546
R3563 VSS.n3037 VSS.n2804 175.546
R3564 VSS.n3030 VSS.n2804 175.546
R3565 VSS.n3030 VSS.n3028 175.546
R3566 VSS.n4331 VSS.n4330 175.546
R3567 VSS.n4330 VSS.n4322 175.546
R3568 VSS.n4326 VSS.n4322 175.546
R3569 VSS.n4326 VSS.n1735 175.546
R3570 VSS.n4639 VSS.n1735 175.546
R3571 VSS.n4639 VSS.n1733 175.546
R3572 VSS.n4643 VSS.n1733 175.546
R3573 VSS.n4643 VSS.n1730 175.546
R3574 VSS.n4649 VSS.n1730 175.546
R3575 VSS.n4649 VSS.n1731 175.546
R3576 VSS.n4365 VSS.n4364 175.546
R3577 VSS.n4364 VSS.n2001 175.546
R3578 VSS.n4360 VSS.n2001 175.546
R3579 VSS.n4360 VSS.n2004 175.546
R3580 VSS.n2026 VSS.n2004 175.546
R3581 VSS.n4349 VSS.n2026 175.546
R3582 VSS.n4349 VSS.n2027 175.546
R3583 VSS.n4345 VSS.n2027 175.546
R3584 VSS.n4345 VSS.n2030 175.546
R3585 VSS.n4338 VSS.n2030 175.546
R3586 VSS.n4338 VSS.n2054 175.546
R3587 VSS.n4636 VSS.n1756 175.546
R3588 VSS.n4465 VSS.n1756 175.546
R3589 VSS.n4465 VSS.n4463 175.546
R3590 VSS.n4470 VSS.n4463 175.546
R3591 VSS.n4470 VSS.n4464 175.546
R3592 VSS.n4464 VSS.n4457 175.546
R3593 VSS.n4483 VSS.n4457 175.546
R3594 VSS.n4483 VSS.n4455 175.546
R3595 VSS.n4488 VSS.n4455 175.546
R3596 VSS.n4488 VSS.n4366 175.546
R3597 VSS.n4494 VSS.n4366 175.546
R3598 VSS.n4309 VSS.n4308 169.925
R3599 VSS.n1463 VSS.n1462 163.333
R3600 VSS.n3800 VSS.n3799 163.333
R3601 VSS.n1563 VSS.n1562 163.333
R3602 VSS.n1584 VSS.n1583 163.333
R3603 VSS.n1171 VSS.n1170 163.333
R3604 VSS.n3606 VSS.n3602 163.333
R3605 VSS.n1408 VSS.n1228 152.643
R3606 VSS.t71 VSS.t28 151.338
R3607 VSS.n1897 VSS.n1896 150
R3608 VSS.n1939 VSS.n1938 150
R3609 VSS.n1909 VSS.n1908 150
R3610 VSS.n1925 VSS.n1257 150
R3611 VSS.n4776 VSS.n1256 150
R3612 VSS.n1452 VSS.n1451 150
R3613 VSS.n1456 VSS.n1455 150
R3614 VSS.n1460 VSS.n1459 150
R3615 VSS.n4773 VSS.n1275 150
R3616 VSS.n1420 VSS.n1419 150
R3617 VSS.n1435 VSS.n1434 150
R3618 VSS.n1443 VSS.n1442 150
R3619 VSS.n4725 VSS.n4724 150
R3620 VSS.n4729 VSS.n4728 150
R3621 VSS.n4733 VSS.n4732 150
R3622 VSS.n4735 VSS.n1274 150
R3623 VSS.n4715 VSS.n1642 150
R3624 VSS.n4715 VSS.n1643 150
R3625 VSS.n1794 VSS.n1793 150
R3626 VSS.n1805 VSS.n1804 150
R3627 VSS.n1814 VSS.n1627 150
R3628 VSS.n4706 VSS.n4705 150
R3629 VSS.n4702 VSS.n4701 150
R3630 VSS.n4698 VSS.n4697 150
R3631 VSS.n4694 VSS.n4693 150
R3632 VSS.n1899 VSS.n1624 150
R3633 VSS.n1935 VSS.n1934 150
R3634 VSS.n1913 VSS.n1912 150
R3635 VSS.n1923 VSS.n1922 150
R3636 VSS.n1722 VSS.n1721 150
R3637 VSS.n1718 VSS.n1717 150
R3638 VSS.n1714 VSS.n1713 150
R3639 VSS.n1710 VSS.n1709 150
R3640 VSS.n4357 VSS.n4356 150
R3641 VSS.n4353 VSS.n4352 150
R3642 VSS.n2033 VSS.n2032 150
R3643 VSS.n4342 VSS.n1650 150
R3644 VSS.n2049 VSS.n2048 150
R3645 VSS.n2045 VSS.n2044 150
R3646 VSS.n2041 VSS.n2040 150
R3647 VSS.n2037 VSS.n2036 150
R3648 VSS.n4712 VSS.n1646 150
R3649 VSS.n4712 VSS.n1647 150
R3650 VSS.n1800 VSS.n1799 150
R3651 VSS.n1811 VSS.n1810 150
R3652 VSS.n1820 VSS.n1819 150
R3653 VSS.n2016 VSS.n2015 150
R3654 VSS.n2012 VSS.n2011 150
R3655 VSS.n2008 VSS.n2007 150
R3656 VSS.n4710 VSS.n1665 150
R3657 VSS.n4459 VSS.n1761 150
R3658 VSS.n4474 VSS.n4473 150
R3659 VSS.n4480 VSS.n4479 150
R3660 VSS.n4453 VSS.n1765 150
R3661 VSS.n4449 VSS.n4448 150
R3662 VSS.n4445 VSS.n4444 150
R3663 VSS.n4441 VSS.n4440 150
R3664 VSS.n4437 VSS.n4436 150
R3665 VSS.n4628 VSS.n1762 150
R3666 VSS.n1828 VSS.n1762 150
R3667 VSS.n4410 VSS.n4409 150
R3668 VSS.n4419 VSS.n4418 150
R3669 VSS.n4428 VSS.n4427 150
R3670 VSS.n2910 VSS.n2909 150
R3671 VSS.n2914 VSS.n2913 150
R3672 VSS.n2918 VSS.n2917 150
R3673 VSS.n2920 VSS.n1779 150
R3674 VSS.n3049 VSS.n3048 150
R3675 VSS.n3045 VSS.n3044 150
R3676 VSS.n2807 VSS.n2806 150
R3677 VSS.n3034 VSS.n2403 150
R3678 VSS.n2822 VSS.n2821 150
R3679 VSS.n2826 VSS.n2825 150
R3680 VSS.n2830 VSS.n2829 150
R3681 VSS.n2834 VSS.n2833 150
R3682 VSS.n3430 VSS.n3429 150
R3683 VSS.n3429 VSS.n2398 150
R3684 VSS.n2878 VSS.n2877 150
R3685 VSS.n2887 VSS.n2886 150
R3686 VSS.n2896 VSS.n2895 150
R3687 VSS.n2790 VSS.n2789 150
R3688 VSS.n2786 VSS.n2785 150
R3689 VSS.n3427 VSS.n2418 150
R3690 VSS.n3423 VSS.n2417 150
R3691 VSS.n2719 VSS.n2718 150
R3692 VSS.n3080 VSS.n3079 150
R3693 VSS.n2728 VSS.n2727 150
R3694 VSS.n3069 VSS.n2472 150
R3695 VSS.n2742 VSS.n2741 150
R3696 VSS.n2738 VSS.n2737 150
R3697 VSS.n2734 VSS.n2733 150
R3698 VSS.n2730 VSS.n2468 150
R3699 VSS.n3375 VSS.n2469 150
R3700 VSS.n2490 VSS.n2469 150
R3701 VSS.n3251 VSS.n3250 150
R3702 VSS.n3260 VSS.n3259 150
R3703 VSS.n3378 VSS.n2467 150
R3704 VSS.n2710 VSS.n2709 150
R3705 VSS.n2706 VSS.n2705 150
R3706 VSS.n2702 VSS.n2701 150
R3707 VSS.n2698 VSS.n2486 150
R3708 VSS.n3914 VSS.n2222 150
R3709 VSS.n2360 VSS.n2359 150
R3710 VSS.n2368 VSS.n2367 150
R3711 VSS.n2342 VSS.n2228 150
R3712 VSS.n2437 VSS.n2436 150
R3713 VSS.n2433 VSS.n2432 150
R3714 VSS.n2429 VSS.n2428 150
R3715 VSS.n2425 VSS.n2242 150
R3716 VSS.n3911 VSS.n2225 150
R3717 VSS.n2248 VSS.n2225 150
R3718 VSS.n3481 VSS.n3480 150
R3719 VSS.n3492 VSS.n3491 150
R3720 VSS.n3502 VSS.n3501 150
R3721 VSS.n3451 VSS.n3450 150
R3722 VSS.n3455 VSS.n3454 150
R3723 VSS.n3459 VSS.n3458 150
R3724 VSS.n3463 VSS.n3462 150
R3725 VSS.n3433 VSS.n2392 150
R3726 VSS.n2868 VSS.n2867 150
R3727 VSS.n2860 VSS.n2859 150
R3728 VSS.n2856 VSS.n2855 150
R3729 VSS.n2456 VSS.n2455 150
R3730 VSS.n2452 VSS.n2451 150
R3731 VSS.n2448 VSS.n2447 150
R3732 VSS.n2444 VSS.n2443 150
R3733 VSS.n2385 VSS.n2384 150
R3734 VSS.n2350 VSS.n2349 150
R3735 VSS.n2347 VSS.n2340 150
R3736 VSS.n2377 VSS.n2333 150
R3737 VSS.n3435 VSS.n2333 150
R3738 VSS.n2848 VSS.n2847 150
R3739 VSS.n2844 VSS.n2843 150
R3740 VSS.n2840 VSS.n2839 150
R3741 VSS.n2836 VSS.n2334 150
R3742 VSS.n5436 VSS.n100 150
R3743 VSS.n5404 VSS.n5403 150
R3744 VSS.n142 VSS.n141 150
R3745 VSS.n5391 VSS.n5390 150
R3746 VSS.n4176 VSS.n4175 150
R3747 VSS.n4180 VSS.n4179 150
R3748 VSS.n4184 VSS.n4183 150
R3749 VSS.n4188 VSS.n4187 150
R3750 VSS.n5453 VSS.n5452 150
R3751 VSS.n85 VSS.n84 150
R3752 VSS.n5438 VSS.n79 150
R3753 VSS.n89 VSS.n80 150
R3754 VSS.n542 VSS.n89 150
R3755 VSS.n443 VSS.n442 150
R3756 VSS.n447 VSS.n446 150
R3757 VSS.n451 VSS.n450 150
R3758 VSS.n455 VSS.n454 150
R3759 VSS.n35 VSS.n34 150
R3760 VSS.n5463 VSS.n37 150
R3761 VSS.n5461 VSS.n38 150
R3762 VSS.n516 VSS.n473 150
R3763 VSS.n5483 VSS.n17 150
R3764 VSS.n5487 VSS.n5485 150
R3765 VSS.n5491 VSS.n15 150
R3766 VSS.n5495 VSS.n5493 150
R3767 VSS.n5506 VSS.n9 150
R3768 VSS.n5508 VSS.n5506 150
R3769 VSS.n5516 VSS.n3 150
R3770 VSS.n5518 VSS.n2 150
R3771 VSS.n499 VSS.n481 150
R3772 VSS.n513 VSS.n474 150
R3773 VSS.n509 VSS.n508 150
R3774 VSS.n506 VSS.n477 150
R3775 VSS.n502 VSS.n501 150
R3776 VSS.n5456 VSS.n61 150
R3777 VSS.n74 VSS.n73 150
R3778 VSS.n5442 VSS.n5441 150
R3779 VSS.n555 VSS.n554 150
R3780 VSS.n4171 VSS.n4170 150
R3781 VSS.n4167 VSS.n4166 150
R3782 VSS.n4163 VSS.n4162 150
R3783 VSS.n4159 VSS.n4158 150
R3784 VSS.n5474 VSS.n5473 150
R3785 VSS.n46 VSS.n45 150
R3786 VSS.n5458 VSS.n40 150
R3787 VSS.n50 VSS.n41 150
R3788 VSS.n458 VSS.n50 150
R3789 VSS.n539 VSS.n538 150
R3790 VSS.n535 VSS.n534 150
R3791 VSS.n531 VSS.n530 150
R3792 VSS.n527 VSS.n526 150
R3793 VSS.n5169 VSS.n5167 150
R3794 VSS.n3687 VSS.n3685 150
R3795 VSS.n3708 VSS.n3674 150
R3796 VSS.n3729 VSS.n3710 150
R3797 VSS.n3726 VSS.n3712 150
R3798 VSS.n3722 VSS.n3721 150
R3799 VSS.n3719 VSS.n3716 150
R3800 VSS.n5228 VSS.n317 150
R3801 VSS.n5197 VSS.n325 150
R3802 VSS.n5208 VSS.n325 150
R3803 VSS.n5212 VSS.n5210 150
R3804 VSS.n5223 VSS.n320 150
R3805 VSS.n5226 VSS.n5225 150
R3806 VSS.n5182 VSS.n5180 150
R3807 VSS.n5186 VSS.n333 150
R3808 VSS.n5190 VSS.n5188 150
R3809 VSS.n5195 VSS.n331 150
R3810 VSS.n370 VSS.n363 150
R3811 VSS.n5149 VSS.n5148 150
R3812 VSS.n3764 VSS.n3763 150
R3813 VSS.n3773 VSS.n3772 150
R3814 VSS.n3784 VSS.n3783 150
R3815 VSS.n3788 VSS.n3787 150
R3816 VSS.n3792 VSS.n3791 150
R3817 VSS.n3796 VSS.n3795 150
R3818 VSS.n357 VSS.n345 150
R3819 VSS.n5164 VSS.n344 150
R3820 VSS.n3691 VSS.n3690 150
R3821 VSS.n3705 VSS.n3704 150
R3822 VSS.n435 VSS.n434 150
R3823 VSS.n431 VSS.n430 150
R3824 VSS.n427 VSS.n426 150
R3825 VSS.n423 VSS.n422 150
R3826 VSS.n5143 VSS.n396 150
R3827 VSS.n5111 VSS.n5110 150
R3828 VSS.n642 VSS.n641 150
R3829 VSS.n5098 VSS.n5097 150
R3830 VSS.n627 VSS.n626 150
R3831 VSS.n623 VSS.n622 150
R3832 VSS.n619 VSS.n618 150
R3833 VSS.n615 VSS.n614 150
R3834 VSS.n5158 VSS.n5157 150
R3835 VSS.n379 VSS.n378 150
R3836 VSS.n5145 VSS.n377 150
R3837 VSS.n3754 VSS.n385 150
R3838 VSS.n3750 VSS.n385 150
R3839 VSS.n3736 VSS.n3735 150
R3840 VSS.n3740 VSS.n3739 150
R3841 VSS.n3744 VSS.n3743 150
R3842 VSS.n3748 VSS.n3747 150
R3843 VSS.n4823 VSS.n918 150
R3844 VSS.n1351 VSS.n919 150
R3845 VSS.n1349 VSS.n1348 150
R3846 VSS.n1344 VSS.n922 150
R3847 VSS.n1189 VSS.n1188 150
R3848 VSS.n1193 VSS.n1192 150
R3849 VSS.n1197 VSS.n1196 150
R3850 VSS.n1199 VSS.n937 150
R3851 VSS.n4820 VSS.n920 150
R3852 VSS.n4812 VSS.n920 150
R3853 VSS.n4809 VSS.n4808 150
R3854 VSS.n4800 VSS.n4799 150
R3855 VSS.n4796 VSS.n4795 150
R3856 VSS.n1337 VSS.n1336 150
R3857 VSS.n1333 VSS.n1332 150
R3858 VSS.n1329 VSS.n1328 150
R3859 VSS.n1325 VSS.n1324 150
R3860 VSS.n1296 VSS.n893 150
R3861 VSS.n1603 VSS.n1602 150
R3862 VSS.n1309 VSS.n1308 150
R3863 VSS.n1588 VSS.n1587 150
R3864 VSS.n1579 VSS.n1578 150
R3865 VSS.n1575 VSS.n1574 150
R3866 VSS.n1571 VSS.n1570 150
R3867 VSS.n1567 VSS.n1566 150
R3868 VSS.n4831 VSS.n911 150
R3869 VSS.n1358 VSS.n1357 150
R3870 VSS.n1367 VSS.n1366 150
R3871 VSS.n1376 VSS.n1375 150
R3872 VSS.n941 VSS.n940 150
R3873 VSS.n945 VSS.n944 150
R3874 VSS.n949 VSS.n948 150
R3875 VSS.n951 VSS.n910 150
R3876 VSS.n4765 VSS.n1282 150
R3877 VSS.n1413 VSS.n1283 150
R3878 VSS.n1439 VSS.n1438 150
R3879 VSS.n1447 VSS.n1446 150
R3880 VSS.n1478 VSS.n1477 150
R3881 VSS.n1474 VSS.n1473 150
R3882 VSS.n1470 VSS.n1469 150
R3883 VSS.n1466 VSS.n1465 150
R3884 VSS.n1614 VSS.n1613 150
R3885 VSS.n1305 VSS.n1304 150
R3886 VSS.n1599 VSS.n1598 150
R3887 VSS.n1318 VSS.n1317 150
R3888 VSS.n4758 VSS.n4757 150
R3889 VSS.n4754 VSS.n4753 150
R3890 VSS.n4750 VSS.n4749 150
R3891 VSS.n4746 VSS.n4745 150
R3892 VSS.n4960 VSS.n724 150
R3893 VSS.n1069 VSS.n1044 150
R3894 VSS.n1073 VSS.n1071 150
R3895 VSS.n1085 VSS.n1038 150
R3896 VSS.n1099 VSS.n1098 150
R3897 VSS.n1096 VSS.n1087 150
R3898 VSS.n1092 VSS.n1091 150
R3899 VSS.n5320 VSS.n279 150
R3900 VSS.n5289 VSS.n287 150
R3901 VSS.n5300 VSS.n287 150
R3902 VSS.n5304 VSS.n5302 150
R3903 VSS.n5315 VSS.n282 150
R3904 VSS.n5318 VSS.n5317 150
R3905 VSS.n4954 VSS.n4940 150
R3906 VSS.n4950 VSS.n4948 150
R3907 VSS.n4946 VSS.n4943 150
R3908 VSS.n5287 VSS.n291 150
R3909 VSS.n752 VSS.n745 150
R3910 VSS.n4921 VSS.n4920 150
R3911 VSS.n1136 VSS.n1135 150
R3912 VSS.n1145 VSS.n1144 150
R3913 VSS.n1156 VSS.n1155 150
R3914 VSS.n1160 VSS.n1159 150
R3915 VSS.n1164 VSS.n1163 150
R3916 VSS.n1168 VSS.n1167 150
R3917 VSS.n728 VSS.n727 150
R3918 VSS.n1052 VSS.n1051 150
R3919 VSS.n1066 VSS.n1065 150
R3920 VSS.n1076 VSS.n1075 150
R3921 VSS.n817 VSS.n816 150
R3922 VSS.n813 VSS.n812 150
R3923 VSS.n809 VSS.n808 150
R3924 VSS.n4936 VSS.n726 150
R3925 VSS.n4915 VSS.n781 150
R3926 VSS.n4883 VSS.n4882 150
R3927 VSS.n849 VSS.n848 150
R3928 VSS.n4870 VSS.n4869 150
R3929 VSS.n835 VSS.n834 150
R3930 VSS.n831 VSS.n830 150
R3931 VSS.n827 VSS.n826 150
R3932 VSS.n823 VSS.n822 150
R3933 VSS.n4930 VSS.n4929 150
R3934 VSS.n764 VSS.n763 150
R3935 VSS.n4917 VSS.n762 150
R3936 VSS.n1126 VSS.n770 150
R3937 VSS.n1122 VSS.n770 150
R3938 VSS.n1108 VSS.n1107 150
R3939 VSS.n1112 VSS.n1111 150
R3940 VSS.n1116 VSS.n1115 150
R3941 VSS.n1120 VSS.n1119 150
R3942 VSS.n3834 VSS.n3832 150
R3943 VSS.n3836 VSS.n3629 150
R3944 VSS.n3611 VSS.n3610 150
R3945 VSS.n3613 VSS.n3609 150
R3946 VSS.n3597 VSS.n3596 150
R3947 VSS.n3594 VSS.n3585 150
R3948 VSS.n3590 VSS.n3589 150
R3949 VSS.n5274 VSS.n298 150
R3950 VSS.n5243 VSS.n306 150
R3951 VSS.n5254 VSS.n306 150
R3952 VSS.n5258 VSS.n5256 150
R3953 VSS.n5269 VSS.n301 150
R3954 VSS.n5272 VSS.n5271 150
R3955 VSS.n3827 VSS.n3813 150
R3956 VSS.n3823 VSS.n3821 150
R3957 VSS.n3819 VSS.n3816 150
R3958 VSS.n5241 VSS.n310 150
R3959 VSS.n3869 VSS.n3867 150
R3960 VSS.n3871 VSS.n2265 150
R3961 VSS.n3555 VSS.n2314 150
R3962 VSS.n3559 VSS.n3557 150
R3963 VSS.n3570 VSS.n2307 150
R3964 VSS.n3574 VSS.n3572 150
R3965 VSS.n3578 VSS.n2305 150
R3966 VSS.n3581 VSS.n3580 150
R3967 VSS.n3846 VSS.n2274 150
R3968 VSS.n3624 VSS.n3623 150
R3969 VSS.n3626 VSS.n3621 150
R3970 VSS.n3604 VSS.n3603 150
R3971 VSS.n3862 VSS.n2270 150
R3972 VSS.n3858 VSS.n3856 150
R3973 VSS.n3854 VSS.n2272 150
R3974 VSS.n3850 VSS.n3848 150
R3975 VSS.n3901 VSS.n3900 150
R3976 VSS.n3903 VSS.n2250 150
R3977 VSS.n3495 VSS.n3470 150
R3978 VSS.n3499 VSS.n3497 150
R3979 VSS.n3897 VSS.n2252 150
R3980 VSS.n3893 VSS.n3891 150
R3981 VSS.n3889 VSS.n2254 150
R3982 VSS.n3885 VSS.n3883 150
R3983 VSS.n3881 VSS.n2256 150
R3984 VSS.n3534 VSS.n3533 150
R3985 VSS.n3550 VSS.n3536 150
R3986 VSS.n3552 VSS.n3531 150
R3987 VSS.n3531 VSS.n3530 150
R3988 VSS.n3517 VSS.n3515 150
R3989 VSS.n3521 VSS.n2319 150
R3990 VSS.n3524 VSS.n3523 150
R3991 VSS.n3528 VSS.n3527 150
R3992 VSS.n3991 VSS.n3990 150
R3993 VSS.n2128 VSS.n2127 150
R3994 VSS.n3978 VSS.n3977 150
R3995 VSS.n2140 VSS.n109 150
R3996 VSS.n5430 VSS.n124 150
R3997 VSS.n5426 VSS.n5425 150
R3998 VSS.n5422 VSS.n5421 150
R3999 VSS.n5418 VSS.n5417 150
R4000 VSS.n5433 VSS.n5432 150
R4001 VSS.n5432 VSS.n104 150
R4002 VSS.n5400 VSS.n5399 150
R4003 VSS.n146 VSS.n145 150
R4004 VSS.n5387 VSS.n5386 150
R4005 VSS.n2165 VSS.n2164 150
R4006 VSS.n2161 VSS.n2160 150
R4007 VSS.n2157 VSS.n2156 150
R4008 VSS.n2153 VSS.n2152 150
R4009 VSS.n4005 VSS.n2085 150
R4010 VSS.n2542 VSS.n2541 150
R4011 VSS.n2568 VSS.n2567 150
R4012 VSS.n2554 VSS.n2553 150
R4013 VSS.n2107 VSS.n2106 150
R4014 VSS.n2111 VSS.n2110 150
R4015 VSS.n4003 VSS.n2104 150
R4016 VSS.n3999 VSS.n2103 150
R4017 VSS.n2122 VSS.n2121 150
R4018 VSS.n3987 VSS.n3986 150
R4019 VSS.n2137 VSS.n2136 150
R4020 VSS.n3974 VSS.n2093 150
R4021 VSS.n2148 VSS.n2093 150
R4022 VSS.n2512 VSS.n2511 150
R4023 VSS.n2508 VSS.n2507 150
R4024 VSS.n2504 VSS.n2503 150
R4025 VSS.n2500 VSS.n2499 150
R4026 VSS.n3211 VSS.n3210 150
R4027 VSS.n3335 VSS.n3334 150
R4028 VSS.n3219 VSS.n3218 150
R4029 VSS.n3318 VSS.n405 150
R4030 VSS.n5137 VSS.n420 150
R4031 VSS.n5133 VSS.n5132 150
R4032 VSS.n5129 VSS.n5128 150
R4033 VSS.n5125 VSS.n5124 150
R4034 VSS.n5140 VSS.n5139 150
R4035 VSS.n5139 VSS.n400 150
R4036 VSS.n5107 VSS.n5106 150
R4037 VSS.n646 VSS.n645 150
R4038 VSS.n5094 VSS.n5093 150
R4039 VSS.n3304 VSS.n3303 150
R4040 VSS.n3300 VSS.n3299 150
R4041 VSS.n3296 VSS.n3295 150
R4042 VSS.n3292 VSS.n3291 150
R4043 VSS.n3365 VSS.n3364 150
R4044 VSS.n3367 VSS.n2492 150
R4045 VSS.n3241 VSS.n3239 150
R4046 VSS.n3269 VSS.n3235 150
R4047 VSS.n3361 VSS.n3195 150
R4048 VSS.n3357 VSS.n3355 150
R4049 VSS.n3353 VSS.n3197 150
R4050 VSS.n3349 VSS.n3347 150
R4051 VSS.n3345 VSS.n3199 150
R4052 VSS.n3329 VSS.n3328 150
R4053 VSS.n3331 VSS.n3326 150
R4054 VSS.n3316 VSS.n3229 150
R4055 VSS.n3316 VSS.n3315 150
R4056 VSS.n3277 VSS.n3274 150
R4057 VSS.n3281 VSS.n3279 150
R4058 VSS.n3285 VSS.n3233 150
R4059 VSS.n3288 VSS.n3287 150
R4060 VSS.n1847 VSS.n1846 150
R4061 VSS.n4588 VSS.n4587 150
R4062 VSS.n1855 VSS.n1854 150
R4063 VSS.n4571 VSS.n790 150
R4064 VSS.n4909 VSS.n805 150
R4065 VSS.n4905 VSS.n4904 150
R4066 VSS.n4901 VSS.n4900 150
R4067 VSS.n4897 VSS.n4896 150
R4068 VSS.n4912 VSS.n4911 150
R4069 VSS.n4911 VSS.n785 150
R4070 VSS.n4879 VSS.n4878 150
R4071 VSS.n853 VSS.n852 150
R4072 VSS.n4866 VSS.n4865 150
R4073 VSS.n1882 VSS.n1881 150
R4074 VSS.n1878 VSS.n1877 150
R4075 VSS.n1874 VSS.n1873 150
R4076 VSS.n1870 VSS.n1869 150
R4077 VSS.n4618 VSS.n4617 150
R4078 VSS.n4620 VSS.n1830 150
R4079 VSS.n4400 VSS.n4398 150
R4080 VSS.n4396 VSS.n4395 150
R4081 VSS.n4614 VSS.n1832 150
R4082 VSS.n4610 VSS.n4608 150
R4083 VSS.n4606 VSS.n1834 150
R4084 VSS.n4602 VSS.n4600 150
R4085 VSS.n4598 VSS.n1836 150
R4086 VSS.n4582 VSS.n4581 150
R4087 VSS.n4584 VSS.n4579 150
R4088 VSS.n4569 VSS.n1865 150
R4089 VSS.n4569 VSS.n4568 150
R4090 VSS.n4390 VSS.n4372 150
R4091 VSS.n4386 VSS.n4385 150
R4092 VSS.n4383 VSS.n4375 150
R4093 VSS.n4379 VSS.n4378 150
R4094 VSS.n2632 VSS.n2631 150
R4095 VSS.n3115 VSS.n3114 150
R4096 VSS.n2641 VSS.n2640 150
R4097 VSS.n3104 VSS.n2524 150
R4098 VSS.n2655 VSS.n2654 150
R4099 VSS.n2651 VSS.n2650 150
R4100 VSS.n2647 VSS.n2646 150
R4101 VSS.n2643 VSS.n2520 150
R4102 VSS.n3143 VSS.n2521 150
R4103 VSS.n2576 VSS.n2521 150
R4104 VSS.n2545 VSS.n2532 150
R4105 VSS.n2564 VSS.n2563 150
R4106 VSS.n3146 VSS.n2519 150
R4107 VSS.n3130 VSS.n3129 150
R4108 VSS.n3134 VSS.n3133 150
R4109 VSS.n3138 VSS.n3137 150
R4110 VSS.n3142 VSS.n3141 150
R4111 VSS.n4305 VSS.n4304 147.656
R4112 VSS.n4276 VSS.n4274 147.339
R4113 VSS.n4261 VSS.n4258 145.082
R4114 VSS.n4258 VSS.n4253 144.706
R4115 VSS.t10 VSS.t6 136.799
R4116 VSS.n1486 VSS.n1226 132.721
R4117 VSS.n4276 VSS.n4275 131.463
R4118 VSS.n5016 VSS.n700 130.291
R4119 VSS.n986 VSS.n960 130.291
R4120 VSS.n1984 VSS.n1956 130.291
R4121 VSS.n2988 VSS.n2966 130.291
R4122 VSS.n597 VSS.n576 130.291
R4123 VSS.n261 VSS.n241 130.291
R4124 VSS.n3635 VSS.n3634 130.291
R4125 VSS.n4995 VSS.n4976 130.291
R4126 VSS.n999 VSS.t32 129.871
R4127 VSS.n218 VSS.t32 129.871
R4128 VSS.n5377 VSS.t32 129.871
R4129 VSS.n5084 VSS.t32 129.871
R4130 VSS.n5047 VSS.t32 129.871
R4131 VSS.n4856 VSS.t32 129.871
R4132 VSS.n2205 VSS.t32 129.871
R4133 VSS.n3923 VSS.t32 129.871
R4134 VSS.n2931 VSS.t32 129.871
R4135 VSS.n4559 VSS.t32 129.871
R4136 VSS.n3418 VSS.t32 129.871
R4137 VSS.t35 VSS.n1745 129.871
R4138 VSS.t35 VSS.n1748 129.871
R4139 VSS.t35 VSS.n1744 129.871
R4140 VSS.n998 VSS.t32 129
R4141 VSS.n5350 VSS.t32 129
R4142 VSS.n5367 VSS.t32 129
R4143 VSS.n5074 VSS.t32 129
R4144 VSS.n5037 VSS.t32 129
R4145 VSS.n4846 VSS.t32 129
R4146 VSS.n2197 VSS.t32 129
R4147 VSS.n3922 VSS.t32 129
R4148 VSS.n2930 VSS.t32 129
R4149 VSS.n4551 VSS.t32 129
R4150 VSS.n3415 VSS.t32 129
R4151 VSS.t35 VSS.n1749 129
R4152 VSS.t35 VSS.n1743 129
R4153 VSS.t35 VSS.n1752 129
R4154 VSS.n5026 VSS.n700 128.599
R4155 VSS.n995 VSS.n960 128.599
R4156 VSS.n4525 VSS.n1956 128.599
R4157 VSS.n2998 VSS.n2966 128.599
R4158 VSS.n607 VSS.n576 128.599
R4159 VSS.n5333 VSS.n241 128.599
R4160 VSS.n3636 VSS.n3635 128.599
R4161 VSS.n5005 VSS.n4976 128.599
R4162 VSS.n4280 VSS.n4268 125.365
R4163 VSS.n1536 VSS.n1382 124.832
R4164 VSS.n4782 VSS.n1249 124.832
R4165 VSS.n4037 VSS.n2066 124.832
R4166 VSS.t89 VSS.t73 120.151
R4167 VSS.t20 VSS.t75 120.093
R4168 VSS.t22 VSS.t8 120.093
R4169 VSS.t2 VSS.t38 118.373
R4170 VSS.t0 VSS.t2 118.373
R4171 VSS.t4 VSS.t0 118.373
R4172 VSS.t28 VSS.t4 118.373
R4173 VSS.n4290 VSS.n4289 117.469
R4174 VSS.n4287 VSS.n4286 116.493
R4175 VSS.n4243 VSS.n4242 116.469
R4176 VSS.n4242 VSS.n4240 112.596
R4177 VSS.t72 VSS.t87 112.138
R4178 VSS.t7 VSS.t9 109.294
R4179 VSS.t68 VSS.t12 109.294
R4180 VSS.t80 VSS.n4237 107.124
R4181 VSS.n4290 VSS.n4239 106.951
R4182 VSS.n4296 VSS.t71 106.385
R4183 VSS.n1408 VSS.n1227 105.951
R4184 VSS.n4297 VSS.t30 105.88
R4185 VSS.n3097 VSS.n2661 103.938
R4186 VSS.t16 VSS.n4257 103.454
R4187 VSS.n5361 VSS.n182 98.5005
R4188 VSS.n5359 VSS.n189 98.5005
R4189 VSS.n693 VSS.n188 98.5005
R4190 VSS.n886 VSS.n187 98.5005
R4191 VSS.n1511 VSS.n1386 98.5005
R4192 VSS.n5340 VSS.n228 98.5005
R4193 VSS.n3805 VSS.n221 98.5005
R4194 VSS.n718 VSS.n227 98.5005
R4195 VSS.n1177 VSS.n226 98.5005
R4196 VSS.n1557 VSS.n1536 98.5005
R4197 VSS.n5381 VSS.n156 98.5005
R4198 VSS.n5088 VSS.n656 98.5005
R4199 VSS.n5050 VSS.n668 98.5005
R4200 VSS.n4860 VSS.n667 98.5005
R4201 VSS.n1485 VSS.n1484 98.5005
R4202 VSS.n3963 VSS.n3962 98.5005
R4203 VSS.n3960 VSS.n2214 98.5005
R4204 VSS.n3443 VSS.n2213 98.5005
R4205 VSS.n4563 VSS.n1890 98.5005
R4206 VSS.n4782 VSS.n1250 98.5005
R4207 VSS.n3153 VSS.n1703 98.5005
R4208 VSS.n3385 VSS.n1704 98.5005
R4209 VSS.n2904 VSS.n1705 98.5005
R4210 VSS.n1964 VSS.n1706 98.5005
R4211 VSS.n4686 VSS.n1708 98.5005
R4212 VSS.n700 VSS.t32 98.0409
R4213 VSS.n960 VSS.t32 98.0409
R4214 VSS.n1956 VSS.t32 98.0409
R4215 VSS.n2966 VSS.t32 98.0409
R4216 VSS.n576 VSS.t32 98.0409
R4217 VSS.n241 VSS.t32 98.0409
R4218 VSS.n3635 VSS.t32 98.0409
R4219 VSS.n4976 VSS.t32 98.0409
R4220 VSS.n2663 VSS.n2660 97.5252
R4221 VSS.n494 VSS.n269 97.5252
R4222 VSS.n5235 VSS.n5234 97.5252
R4223 VSS.n5327 VSS.n5326 97.5252
R4224 VSS.n5281 VSS.n5280 97.5252
R4225 VSS.n3063 VSS.n2747 97.5252
R4226 VSS.n3028 VSS.n1755 97.5252
R4227 VSS.n4495 VSS.n4494 97.5252
R4228 VSS.t26 VSS.t66 96.2189
R4229 VSS.t11 VSS.t86 94.772
R4230 VSS.n4199 VSS.n4197 93.6243
R4231 VSS.n572 VSS.n180 93.6243
R4232 VSS.n5356 VSS.n184 93.6243
R4233 VSS.n5030 VSS.n185 93.6243
R4234 VSS.n4839 VSS.n186 93.6243
R4235 VSS.n4135 VSS.n4097 93.6243
R4236 VSS.n5337 VSS.n223 93.6243
R4237 VSS.n5342 VSS.n222 93.6243
R4238 VSS.n5009 VSS.n224 93.6243
R4239 VSS.n1179 VSS.n225 93.6243
R4240 VSS.n5413 VSS.n128 93.6243
R4241 VSS.n5120 VSS.n630 93.6243
R4242 VSS.n5052 VSS.n663 93.6243
R4243 VSS.n4892 VSS.n664 93.6243
R4244 VSS.n4739 VSS.n665 93.6243
R4245 VSS.n4037 VSS.n2067 93.6243
R4246 VSS.n2209 VSS.n2171 93.6243
R4247 VSS.n3957 VSS.n2210 93.6243
R4248 VSS.n2329 VSS.n2211 93.6243
R4249 VSS.n1952 VSS.n1950 93.6243
R4250 VSS.n2600 VSS.n1701 93.6243
R4251 VSS.n2497 VSS.n1695 93.6243
R4252 VSS.n2462 VSS.n1689 93.6243
R4253 VSS.n2928 VSS.n1683 93.6243
R4254 VSS.n4522 VSS.n1677 93.6243
R4255 VSS.t87 VSS.t21 91.9235
R4256 VSS.n5327 VSS.n274 89.7233
R4257 VSS.n327 VSS.n269 89.7233
R4258 VSS.n5283 VSS.n5281 89.7233
R4259 VSS.n5237 VSS.n5235 89.7233
R4260 VSS.n3095 VSS.n2663 89.7233
R4261 VSS.n3057 VSS.n2747 89.7233
R4262 VSS.n4495 VSS.n4365 89.7233
R4263 VSS.n4636 VSS.n1755 89.7233
R4264 VSS.n5349 VSS.n202 87.7728
R4265 VSS.n3184 VSS.n2495 87.7728
R4266 VSS.n3184 VSS.n3157 87.7728
R4267 VSS.n3180 VSS.n3157 87.7728
R4268 VSS.n3180 VSS.n3177 87.7728
R4269 VSS.n3177 VSS.n3176 87.7728
R4270 VSS.n3176 VSS.n3159 87.7728
R4271 VSS.n3172 VSS.n3159 87.7728
R4272 VSS.n3172 VSS.n3162 87.7728
R4273 VSS.n3164 VSS.n3162 87.7728
R4274 VSS.n3167 VSS.n3164 87.7728
R4275 VSS.n2692 VSS.n2666 87.7728
R4276 VSS.n2688 VSS.n2666 87.7728
R4277 VSS.n2688 VSS.n2668 87.7728
R4278 VSS.n2684 VSS.n2668 87.7728
R4279 VSS.n2684 VSS.n2683 87.7728
R4280 VSS.n2683 VSS.n2682 87.7728
R4281 VSS.n2682 VSS.n2671 87.7728
R4282 VSS.n2678 VSS.n2671 87.7728
R4283 VSS.n2678 VSS.n2674 87.7728
R4284 VSS.n2674 VSS.n2496 87.7728
R4285 VSS.n4301 VSS.t39 87.6484
R4286 VSS.t84 VSS.t74 87.5807
R4287 VSS.t85 VSS.t84 81.7903
R4288 VSS.n3060 VSS.n2747 79.9708
R4289 VSS.n3025 VSS.n1755 79.9708
R4290 VSS.n4496 VSS.n4495 79.9708
R4291 VSS.n2696 VSS.n2663 79.9708
R4292 VSS.n4295 VSS.n4293 79.0663
R4293 VSS.n4295 VSS.n4294 78.778
R4294 VSS.t21 VSS.t6 77.4474
R4295 VSS.n1553 VSS.n1240 76.3222
R4296 VSS.n1549 VSS.n1241 76.3222
R4297 VSS.n1545 VSS.n1242 76.3222
R4298 VSS.n1541 VSS.n1243 76.3222
R4299 VSS.n4785 VSS.n1221 76.3222
R4300 VSS.n1512 VSS.n1234 76.3222
R4301 VSS.n1516 VSS.n1235 76.3222
R4302 VSS.n1520 VSS.n1236 76.3222
R4303 VSS.n1524 VSS.n1237 76.3222
R4304 VSS.n1528 VSS.n1238 76.3222
R4305 VSS.n1382 VSS.n1246 76.3222
R4306 VSS.n1491 VSS.n1229 76.3222
R4307 VSS.n1495 VSS.n1230 76.3222
R4308 VSS.n1499 VSS.n1231 76.3222
R4309 VSS.n1503 VSS.n1232 76.3222
R4310 VSS.n1389 VSS.n1222 76.3222
R4311 VSS.n1393 VSS.n1223 76.3222
R4312 VSS.n1397 VSS.n1224 76.3222
R4313 VSS.n1401 VSS.n1225 76.3222
R4314 VSS.n1405 VSS.n1226 76.3222
R4315 VSS.n4652 VSS.n1727 76.3222
R4316 VSS.n4078 VSS.n4076 76.3222
R4317 VSS.n4064 VSS.n4063 76.3222
R4318 VSS.n2599 VSS.n2079 76.3222
R4319 VSS.n4131 VSS.n4092 76.3222
R4320 VSS.n2622 VSS.n2589 76.3222
R4321 VSS.n5500 VSS.n5499 76.3222
R4322 VSS.n5503 VSS.n5502 76.3222
R4323 VSS.n5512 VSS.n5511 76.3222
R4324 VSS.n484 VSS.n5 76.3222
R4325 VSS.n490 VSS.n489 76.3222
R4326 VSS.n496 VSS.n495 76.3222
R4327 VSS.n1206 VSS.n274 76.3222
R4328 VSS.n4817 VSS.n4816 76.3222
R4329 VSS.n1210 VSS.n1208 76.3222
R4330 VSS.n4805 VSS.n4804 76.3222
R4331 VSS.n1216 VSS.n1212 76.3222
R4332 VSS.n4792 VSS.n4791 76.3222
R4333 VSS.n328 VSS.n327 76.3222
R4334 VSS.n5202 VSS.n5201 76.3222
R4335 VSS.n5205 VSS.n5204 76.3222
R4336 VSS.n5217 VSS.n5216 76.3222
R4337 VSS.n5220 VSS.n5219 76.3222
R4338 VSS.n5233 VSS.n5232 76.3222
R4339 VSS.n5283 VSS.n5282 76.3222
R4340 VSS.n5294 VSS.n5293 76.3222
R4341 VSS.n5297 VSS.n5296 76.3222
R4342 VSS.n5309 VSS.n5308 76.3222
R4343 VSS.n5312 VSS.n5311 76.3222
R4344 VSS.n5325 VSS.n5324 76.3222
R4345 VSS.n5237 VSS.n5236 76.3222
R4346 VSS.n5248 VSS.n5247 76.3222
R4347 VSS.n5251 VSS.n5250 76.3222
R4348 VSS.n5263 VSS.n5262 76.3222
R4349 VSS.n5266 VSS.n5265 76.3222
R4350 VSS.n5279 VSS.n5278 76.3222
R4351 VSS.n4332 VSS.n4331 76.3222
R4352 VSS.n5501 VSS.n5500 76.3222
R4353 VSS.n5502 VSS.n7 76.3222
R4354 VSS.n5513 VSS.n5512 76.3222
R4355 VSS.n485 VSS.n484 76.3222
R4356 VSS.n491 VSS.n490 76.3222
R4357 VSS.n495 VSS.n494 76.3222
R4358 VSS.n329 VSS.n328 76.3222
R4359 VSS.n5203 VSS.n5202 76.3222
R4360 VSS.n5204 VSS.n322 76.3222
R4361 VSS.n5218 VSS.n5217 76.3222
R4362 VSS.n5219 VSS.n314 76.3222
R4363 VSS.n5234 VSS.n5233 76.3222
R4364 VSS.n5236 VSS.n308 76.3222
R4365 VSS.n5249 VSS.n5248 76.3222
R4366 VSS.n5250 VSS.n303 76.3222
R4367 VSS.n5264 VSS.n5263 76.3222
R4368 VSS.n5265 VSS.n295 76.3222
R4369 VSS.n5280 VSS.n5279 76.3222
R4370 VSS.n5282 VSS.n289 76.3222
R4371 VSS.n5295 VSS.n5294 76.3222
R4372 VSS.n5296 VSS.n284 76.3222
R4373 VSS.n5310 VSS.n5309 76.3222
R4374 VSS.n5311 VSS.n276 76.3222
R4375 VSS.n5326 VSS.n5325 76.3222
R4376 VSS.n1207 VSS.n1206 76.3222
R4377 VSS.n4816 VSS.n4815 76.3222
R4378 VSS.n1211 VSS.n1210 76.3222
R4379 VSS.n4804 VSS.n4803 76.3222
R4380 VSS.n1217 VSS.n1216 76.3222
R4381 VSS.n4791 VSS.n4790 76.3222
R4382 VSS.n2622 VSS.n2621 76.3222
R4383 VSS.n2079 VSS.n2077 76.3222
R4384 VSS.n4063 VSS.n4061 76.3222
R4385 VSS.n4079 VSS.n4078 76.3222
R4386 VSS.n4131 VSS.n4130 76.3222
R4387 VSS.n4333 VSS.n4332 76.3222
R4388 VSS.n4654 VSS.n1727 76.3222
R4389 VSS.n1404 VSS.n1225 76.3222
R4390 VSS.n1400 VSS.n1224 76.3222
R4391 VSS.n1396 VSS.n1223 76.3222
R4392 VSS.n1392 VSS.n1222 76.3222
R4393 VSS.n1506 VSS.n1232 76.3222
R4394 VSS.n1502 VSS.n1231 76.3222
R4395 VSS.n1498 VSS.n1230 76.3222
R4396 VSS.n1494 VSS.n1229 76.3222
R4397 VSS.n1490 VSS.n1228 76.3222
R4398 VSS.n1532 VSS.n1246 76.3222
R4399 VSS.n1531 VSS.n1238 76.3222
R4400 VSS.n1527 VSS.n1237 76.3222
R4401 VSS.n1523 VSS.n1236 76.3222
R4402 VSS.n1519 VSS.n1235 76.3222
R4403 VSS.n1515 VSS.n1234 76.3222
R4404 VSS.n4786 VSS.n4785 76.3222
R4405 VSS.n1538 VSS.n1243 76.3222
R4406 VSS.n1542 VSS.n1242 76.3222
R4407 VSS.n1546 VSS.n1241 76.3222
R4408 VSS.n1550 VSS.n1240 76.3222
R4409 VSS.n4706 VSS.n1637 76.062
R4410 VSS.n1642 VSS.n1637 76.062
R4411 VSS.n4775 VSS.n1257 74.5978
R4412 VSS.n3773 VSS.n353 74.5978
R4413 VSS.n3783 VSS.n353 74.5978
R4414 VSS.n1588 VSS.n900 74.5978
R4415 VSS.n1447 VSS.n1292 74.5978
R4416 VSS.n1579 VSS.n900 74.5978
R4417 VSS.n1145 VSS.n737 74.5978
R4418 VSS.n1155 VSS.n737 74.5978
R4419 VSS.n3559 VSS.n3558 74.5978
R4420 VSS.n3558 VSS.n2307 74.5978
R4421 VSS.n4776 VSS.n4775 74.5978
R4422 VSS.n1478 VSS.n1292 74.5978
R4423 VSS.t86 VSS.t15 74.5155
R4424 VSS.t66 VSS.t19 73.0686
R4425 VSS.n4286 VSS.n4247 72.0167
R4426 VSS.n4774 VSS.n4773 69.3109
R4427 VSS.n4711 VSS.n1646 69.3109
R4428 VSS.n4711 VSS.n4710 69.3109
R4429 VSS.n4629 VSS.n4628 69.3109
R4430 VSS.n4629 VSS.n1779 69.3109
R4431 VSS.n3430 VSS.n2397 69.3109
R4432 VSS.n3423 VSS.n2397 69.3109
R4433 VSS.n3376 VSS.n3375 69.3109
R4434 VSS.n3376 VSS.n2486 69.3109
R4435 VSS.n3912 VSS.n3911 69.3109
R4436 VSS.n3912 VSS.n2242 69.3109
R4437 VSS.n2386 VSS.n2385 69.3109
R4438 VSS.n2443 VSS.n2386 69.3109
R4439 VSS.n5453 VSS.n64 69.3109
R4440 VSS.n4188 VSS.n64 69.3109
R4441 VSS.n5494 VSS.n9 69.3109
R4442 VSS.n5495 VSS.n5494 69.3109
R4443 VSS.n5474 VSS.n22 69.3109
R4444 VSS.n4158 VSS.n22 69.3109
R4445 VSS.n5197 VSS.n5196 69.3109
R4446 VSS.n358 VSS.n357 69.3109
R4447 VSS.n422 VSS.n358 69.3109
R4448 VSS.n5196 VSS.n5195 69.3109
R4449 VSS.n5158 VSS.n367 69.3109
R4450 VSS.n614 VSS.n367 69.3109
R4451 VSS.n4821 VSS.n4820 69.3109
R4452 VSS.n4821 VSS.n937 69.3109
R4453 VSS.n4832 VSS.n4831 69.3109
R4454 VSS.n1615 VSS.n1614 69.3109
R4455 VSS.n4745 VSS.n1615 69.3109
R4456 VSS.n4832 VSS.n910 69.3109
R4457 VSS.n5289 VSS.n5288 69.3109
R4458 VSS.n4935 VSS.n727 69.3109
R4459 VSS.n4936 VSS.n4935 69.3109
R4460 VSS.n5288 VSS.n5287 69.3109
R4461 VSS.n4930 VSS.n749 69.3109
R4462 VSS.n822 VSS.n749 69.3109
R4463 VSS.n5243 VSS.n5242 69.3109
R4464 VSS.n3847 VSS.n3846 69.3109
R4465 VSS.n3848 VSS.n3847 69.3109
R4466 VSS.n5242 VSS.n5241 69.3109
R4467 VSS.n3882 VSS.n3881 69.3109
R4468 VSS.n3883 VSS.n3882 69.3109
R4469 VSS.n5433 VSS.n103 69.3109
R4470 VSS.n5417 VSS.n103 69.3109
R4471 VSS.n2121 VSS.n2099 69.3109
R4472 VSS.n3999 VSS.n2099 69.3109
R4473 VSS.n5140 VSS.n399 69.3109
R4474 VSS.n5124 VSS.n399 69.3109
R4475 VSS.n3346 VSS.n3345 69.3109
R4476 VSS.n3347 VSS.n3346 69.3109
R4477 VSS.n4912 VSS.n784 69.3109
R4478 VSS.n4896 VSS.n784 69.3109
R4479 VSS.n4599 VSS.n4598 69.3109
R4480 VSS.n4600 VSS.n4599 69.3109
R4481 VSS.n3144 VSS.n3143 69.3109
R4482 VSS.n3144 VSS.n3142 69.3109
R4483 VSS.n4774 VSS.n1274 69.3109
R4484 VSS.t48 VSS.n1628 65.8183
R4485 VSS.t48 VSS.n1629 65.8183
R4486 VSS.t48 VSS.n1630 65.8183
R4487 VSS.t48 VSS.n1631 65.8183
R4488 VSS.t58 VSS.n1651 65.8183
R4489 VSS.t58 VSS.n1652 65.8183
R4490 VSS.t58 VSS.n1653 65.8183
R4491 VSS.t58 VSS.n1654 65.8183
R4492 VSS.t58 VSS.n1661 65.8183
R4493 VSS.t58 VSS.n1662 65.8183
R4494 VSS.t58 VSS.n1663 65.8183
R4495 VSS.t58 VSS.n1664 65.8183
R4496 VSS.t44 VSS.n1766 65.8183
R4497 VSS.t44 VSS.n1767 65.8183
R4498 VSS.t44 VSS.n1768 65.8183
R4499 VSS.t44 VSS.n1769 65.8183
R4500 VSS.t44 VSS.n1775 65.8183
R4501 VSS.t44 VSS.n1776 65.8183
R4502 VSS.t44 VSS.n1777 65.8183
R4503 VSS.t44 VSS.n1778 65.8183
R4504 VSS.t61 VSS.n2404 65.8183
R4505 VSS.t61 VSS.n2405 65.8183
R4506 VSS.t61 VSS.n2406 65.8183
R4507 VSS.t61 VSS.n2407 65.8183
R4508 VSS.t61 VSS.n2414 65.8183
R4509 VSS.t61 VSS.n2415 65.8183
R4510 VSS.t61 VSS.n2416 65.8183
R4511 VSS.t61 VSS.n3428 65.8183
R4512 VSS.t64 VSS.n2473 65.8183
R4513 VSS.t64 VSS.n2474 65.8183
R4514 VSS.t64 VSS.n2475 65.8183
R4515 VSS.t64 VSS.n2476 65.8183
R4516 VSS.t64 VSS.n2482 65.8183
R4517 VSS.t64 VSS.n2483 65.8183
R4518 VSS.t64 VSS.n2484 65.8183
R4519 VSS.t64 VSS.n2485 65.8183
R4520 VSS.t65 VSS.n2241 65.8183
R4521 VSS.t65 VSS.n2240 65.8183
R4522 VSS.t65 VSS.n2239 65.8183
R4523 VSS.t65 VSS.n2238 65.8183
R4524 VSS.t47 VSS.n2387 65.8183
R4525 VSS.t47 VSS.n2388 65.8183
R4526 VSS.t47 VSS.n2389 65.8183
R4527 VSS.t47 VSS.n2390 65.8183
R4528 VSS.t47 VSS.n2383 65.8183
R4529 VSS.t47 VSS.n2382 65.8183
R4530 VSS.t47 VSS.n2381 65.8183
R4531 VSS.t47 VSS.n2380 65.8183
R4532 VSS.t65 VSS.n2229 65.8183
R4533 VSS.t65 VSS.n2230 65.8183
R4534 VSS.t65 VSS.n2231 65.8183
R4535 VSS.t65 VSS.n2232 65.8183
R4536 VSS.t36 VSS.n95 65.8183
R4537 VSS.t36 VSS.n96 65.8183
R4538 VSS.t36 VSS.n97 65.8183
R4539 VSS.t36 VSS.n98 65.8183
R4540 VSS.t36 VSS.n94 65.8183
R4541 VSS.t36 VSS.n93 65.8183
R4542 VSS.t36 VSS.n92 65.8183
R4543 VSS.t36 VSS.n91 65.8183
R4544 VSS.n5478 VSS.t40 65.8183
R4545 VSS.n5484 VSS.t40 65.8183
R4546 VSS.n5486 VSS.t40 65.8183
R4547 VSS.n5492 VSS.t40 65.8183
R4548 VSS.t62 VSS.n56 65.8183
R4549 VSS.t62 VSS.n57 65.8183
R4550 VSS.t62 VSS.n58 65.8183
R4551 VSS.t62 VSS.n59 65.8183
R4552 VSS.t62 VSS.n55 65.8183
R4553 VSS.t62 VSS.n54 65.8183
R4554 VSS.t62 VSS.n53 65.8183
R4555 VSS.t62 VSS.n52 65.8183
R4556 VSS.n479 VSS.t40 65.8183
R4557 VSS.n507 VSS.t40 65.8183
R4558 VSS.n476 VSS.t40 65.8183
R4559 VSS.n514 VSS.t40 65.8183
R4560 VSS.n472 VSS.t40 65.8183
R4561 VSS.n5462 VSS.t40 65.8183
R4562 VSS.n36 VSS.t40 65.8183
R4563 VSS.n19 VSS.t40 65.8183
R4564 VSS.n5457 VSS.t62 65.8183
R4565 VSS.t62 VSS.n47 65.8183
R4566 VSS.t62 VSS.n23 65.8183
R4567 VSS.t62 VSS.n49 65.8183
R4568 VSS.t62 VSS.n48 65.8183
R4569 VSS.t62 VSS.n43 65.8183
R4570 VSS.t62 VSS.n42 65.8183
R4571 VSS.n5437 VSS.t36 65.8183
R4572 VSS.t36 VSS.n86 65.8183
R4573 VSS.t36 VSS.n65 65.8183
R4574 VSS.n3715 VSS.t50 65.8183
R4575 VSS.n3720 VSS.t50 65.8183
R4576 VSS.n3714 VSS.t50 65.8183
R4577 VSS.n3727 VSS.t50 65.8183
R4578 VSS.t41 VSS.n359 65.8183
R4579 VSS.t41 VSS.n360 65.8183
R4580 VSS.t41 VSS.n361 65.8183
R4581 VSS.t41 VSS.n362 65.8183
R4582 VSS.n5179 VSS.t50 65.8183
R4583 VSS.n5181 VSS.t50 65.8183
R4584 VSS.n5187 VSS.t50 65.8183
R4585 VSS.n5189 VSS.t50 65.8183
R4586 VSS.n3709 VSS.t50 65.8183
R4587 VSS.n3686 VSS.t50 65.8183
R4588 VSS.n341 VSS.t50 65.8183
R4589 VSS.n5168 VSS.t50 65.8183
R4590 VSS.t41 VSS.n348 65.8183
R4591 VSS.t41 VSS.n347 65.8183
R4592 VSS.t41 VSS.n346 65.8183
R4593 VSS.n5163 VSS.t41 65.8183
R4594 VSS.t63 VSS.n391 65.8183
R4595 VSS.t63 VSS.n392 65.8183
R4596 VSS.t63 VSS.n393 65.8183
R4597 VSS.t63 VSS.n394 65.8183
R4598 VSS.t63 VSS.n390 65.8183
R4599 VSS.t63 VSS.n389 65.8183
R4600 VSS.t63 VSS.n388 65.8183
R4601 VSS.t63 VSS.n387 65.8183
R4602 VSS.t41 VSS.n352 65.8183
R4603 VSS.t41 VSS.n351 65.8183
R4604 VSS.t41 VSS.n350 65.8183
R4605 VSS.t41 VSS.n349 65.8183
R4606 VSS.t53 VSS.n936 65.8183
R4607 VSS.t53 VSS.n935 65.8183
R4608 VSS.t53 VSS.n934 65.8183
R4609 VSS.t53 VSS.n933 65.8183
R4610 VSS.t60 VSS.n1616 65.8183
R4611 VSS.t60 VSS.n1617 65.8183
R4612 VSS.t60 VSS.n1618 65.8183
R4613 VSS.t60 VSS.n1619 65.8183
R4614 VSS.t45 VSS.n909 65.8183
R4615 VSS.t45 VSS.n908 65.8183
R4616 VSS.t45 VSS.n907 65.8183
R4617 VSS.t45 VSS.n906 65.8183
R4618 VSS.t45 VSS.n898 65.8183
R4619 VSS.t45 VSS.n905 65.8183
R4620 VSS.t45 VSS.n895 65.8183
R4621 VSS.n4833 VSS.t45 65.8183
R4622 VSS.t60 VSS.n1287 65.8183
R4623 VSS.t60 VSS.n1286 65.8183
R4624 VSS.t60 VSS.n1285 65.8183
R4625 VSS.t60 VSS.n1284 65.8183
R4626 VSS.t45 VSS.n904 65.8183
R4627 VSS.t45 VSS.n903 65.8183
R4628 VSS.t45 VSS.n902 65.8183
R4629 VSS.t45 VSS.n901 65.8183
R4630 VSS.t53 VSS.n923 65.8183
R4631 VSS.t53 VSS.n924 65.8183
R4632 VSS.t53 VSS.n925 65.8183
R4633 VSS.t53 VSS.n926 65.8183
R4634 VSS.t53 VSS.n921 65.8183
R4635 VSS.t53 VSS.n929 65.8183
R4636 VSS.n4822 VSS.t53 65.8183
R4637 VSS.t53 VSS.n932 65.8183
R4638 VSS.t45 VSS.n899 65.8183
R4639 VSS.t45 VSS.n897 65.8183
R4640 VSS.t45 VSS.n896 65.8183
R4641 VSS.t45 VSS.n894 65.8183
R4642 VSS.n1090 VSS.t51 65.8183
R4643 VSS.n1089 VSS.t51 65.8183
R4644 VSS.n1097 VSS.t51 65.8183
R4645 VSS.n1100 VSS.t51 65.8183
R4646 VSS.t42 VSS.n741 65.8183
R4647 VSS.t42 VSS.n742 65.8183
R4648 VSS.t42 VSS.n743 65.8183
R4649 VSS.t42 VSS.n744 65.8183
R4650 VSS.n4955 VSS.t51 65.8183
R4651 VSS.n4949 VSS.t51 65.8183
R4652 VSS.n4947 VSS.t51 65.8183
R4653 VSS.n4942 VSS.t51 65.8183
R4654 VSS.n1072 VSS.t51 65.8183
R4655 VSS.n1070 VSS.t51 65.8183
R4656 VSS.n1043 VSS.t51 65.8183
R4657 VSS.n4959 VSS.t51 65.8183
R4658 VSS.t42 VSS.n732 65.8183
R4659 VSS.t42 VSS.n731 65.8183
R4660 VSS.t42 VSS.n730 65.8183
R4661 VSS.t42 VSS.n729 65.8183
R4662 VSS.t46 VSS.n776 65.8183
R4663 VSS.t46 VSS.n777 65.8183
R4664 VSS.t46 VSS.n778 65.8183
R4665 VSS.t46 VSS.n779 65.8183
R4666 VSS.t46 VSS.n775 65.8183
R4667 VSS.t46 VSS.n774 65.8183
R4668 VSS.t46 VSS.n773 65.8183
R4669 VSS.t46 VSS.n772 65.8183
R4670 VSS.t42 VSS.n736 65.8183
R4671 VSS.t42 VSS.n735 65.8183
R4672 VSS.t42 VSS.n734 65.8183
R4673 VSS.t42 VSS.n733 65.8183
R4674 VSS.t42 VSS.n738 65.8183
R4675 VSS.t42 VSS.n739 65.8183
R4676 VSS.t42 VSS.n740 65.8183
R4677 VSS.t42 VSS.n4934 65.8183
R4678 VSS.t46 VSS.n768 65.8183
R4679 VSS.n4916 VSS.t46 65.8183
R4680 VSS.t46 VSS.n750 65.8183
R4681 VSS.n3588 VSS.t57 65.8183
R4682 VSS.n3587 VSS.t57 65.8183
R4683 VSS.n3595 VSS.t57 65.8183
R4684 VSS.n3584 VSS.t57 65.8183
R4685 VSS.n3863 VSS.t52 65.8183
R4686 VSS.n3857 VSS.t52 65.8183
R4687 VSS.n3855 VSS.t52 65.8183
R4688 VSS.n3849 VSS.t52 65.8183
R4689 VSS.n3828 VSS.t57 65.8183
R4690 VSS.n3822 VSS.t57 65.8183
R4691 VSS.n3820 VSS.t57 65.8183
R4692 VSS.n3815 VSS.t57 65.8183
R4693 VSS.n3612 VSS.t57 65.8183
R4694 VSS.n2283 VSS.t57 65.8183
R4695 VSS.n3835 VSS.t57 65.8183
R4696 VSS.n3831 VSS.t57 65.8183
R4697 VSS.n3605 VSS.t52 65.8183
R4698 VSS.n2285 VSS.t52 65.8183
R4699 VSS.n3625 VSS.t52 65.8183
R4700 VSS.n3622 VSS.t52 65.8183
R4701 VSS.n3898 VSS.t59 65.8183
R4702 VSS.n3892 VSS.t59 65.8183
R4703 VSS.n3890 VSS.t59 65.8183
R4704 VSS.n3884 VSS.t59 65.8183
R4705 VSS.n2317 VSS.t59 65.8183
R4706 VSS.n3522 VSS.t59 65.8183
R4707 VSS.n3516 VSS.t59 65.8183
R4708 VSS.n3514 VSS.t59 65.8183
R4709 VSS.n2303 VSS.t52 65.8183
R4710 VSS.n3579 VSS.t52 65.8183
R4711 VSS.n3573 VSS.t52 65.8183
R4712 VSS.n3571 VSS.t52 65.8183
R4713 VSS.n3556 VSS.t52 65.8183
R4714 VSS.n2313 VSS.t52 65.8183
R4715 VSS.n3870 VSS.t52 65.8183
R4716 VSS.n3866 VSS.t52 65.8183
R4717 VSS.n3551 VSS.t59 65.8183
R4718 VSS.n3535 VSS.t59 65.8183
R4719 VSS.n3532 VSS.t59 65.8183
R4720 VSS.t41 VSS.n354 65.8183
R4721 VSS.t41 VSS.n355 65.8183
R4722 VSS.t41 VSS.n356 65.8183
R4723 VSS.t41 VSS.n5162 65.8183
R4724 VSS.t63 VSS.n383 65.8183
R4725 VSS.n5144 VSS.t63 65.8183
R4726 VSS.t63 VSS.n368 65.8183
R4727 VSS.t31 VSS.n5431 65.8183
R4728 VSS.t31 VSS.n122 65.8183
R4729 VSS.t31 VSS.n121 65.8183
R4730 VSS.t31 VSS.n120 65.8183
R4731 VSS.t54 VSS.n2100 65.8183
R4732 VSS.t54 VSS.n2101 65.8183
R4733 VSS.t54 VSS.n2102 65.8183
R4734 VSS.t54 VSS.n4004 65.8183
R4735 VSS.t54 VSS.n2098 65.8183
R4736 VSS.t54 VSS.n2097 65.8183
R4737 VSS.t54 VSS.n2096 65.8183
R4738 VSS.t54 VSS.n2095 65.8183
R4739 VSS.t31 VSS.n110 65.8183
R4740 VSS.t31 VSS.n111 65.8183
R4741 VSS.t31 VSS.n112 65.8183
R4742 VSS.t31 VSS.n113 65.8183
R4743 VSS.t56 VSS.n5138 65.8183
R4744 VSS.t56 VSS.n418 65.8183
R4745 VSS.t56 VSS.n417 65.8183
R4746 VSS.t56 VSS.n416 65.8183
R4747 VSS.n3362 VSS.t49 65.8183
R4748 VSS.n3356 VSS.t49 65.8183
R4749 VSS.n3354 VSS.t49 65.8183
R4750 VSS.n3348 VSS.t49 65.8183
R4751 VSS.n3286 VSS.t49 65.8183
R4752 VSS.n3280 VSS.t49 65.8183
R4753 VSS.n3278 VSS.t49 65.8183
R4754 VSS.n3273 VSS.t49 65.8183
R4755 VSS.t56 VSS.n406 65.8183
R4756 VSS.t56 VSS.n407 65.8183
R4757 VSS.t56 VSS.n408 65.8183
R4758 VSS.t56 VSS.n409 65.8183
R4759 VSS.t56 VSS.n404 65.8183
R4760 VSS.t56 VSS.n412 65.8183
R4761 VSS.t56 VSS.n403 65.8183
R4762 VSS.t56 VSS.n415 65.8183
R4763 VSS.n3216 VSS.t49 65.8183
R4764 VSS.n3330 VSS.t49 65.8183
R4765 VSS.n3327 VSS.t49 65.8183
R4766 VSS.t31 VSS.n108 65.8183
R4767 VSS.t31 VSS.n116 65.8183
R4768 VSS.t31 VSS.n107 65.8183
R4769 VSS.t31 VSS.n119 65.8183
R4770 VSS.t54 VSS.n2091 65.8183
R4771 VSS.t54 VSS.n2089 65.8183
R4772 VSS.t54 VSS.n2087 65.8183
R4773 VSS.t43 VSS.n4910 65.8183
R4774 VSS.t43 VSS.n803 65.8183
R4775 VSS.t43 VSS.n802 65.8183
R4776 VSS.t43 VSS.n801 65.8183
R4777 VSS.n4615 VSS.t33 65.8183
R4778 VSS.n4609 VSS.t33 65.8183
R4779 VSS.n4607 VSS.t33 65.8183
R4780 VSS.n4601 VSS.t33 65.8183
R4781 VSS.n4377 VSS.t33 65.8183
R4782 VSS.n4384 VSS.t33 65.8183
R4783 VSS.n4374 VSS.t33 65.8183
R4784 VSS.n4391 VSS.t33 65.8183
R4785 VSS.t43 VSS.n791 65.8183
R4786 VSS.t43 VSS.n792 65.8183
R4787 VSS.t43 VSS.n793 65.8183
R4788 VSS.t43 VSS.n794 65.8183
R4789 VSS.t43 VSS.n789 65.8183
R4790 VSS.t43 VSS.n797 65.8183
R4791 VSS.t43 VSS.n788 65.8183
R4792 VSS.t43 VSS.n800 65.8183
R4793 VSS.n1852 VSS.t33 65.8183
R4794 VSS.n4583 VSS.t33 65.8183
R4795 VSS.n4580 VSS.t33 65.8183
R4796 VSS.t65 VSS.n2227 65.8183
R4797 VSS.t65 VSS.n2235 65.8183
R4798 VSS.t65 VSS.n2226 65.8183
R4799 VSS.n3913 VSS.t65 65.8183
R4800 VSS.t47 VSS.n2378 65.8183
R4801 VSS.t47 VSS.n2338 65.8183
R4802 VSS.t47 VSS.n2336 65.8183
R4803 VSS.t34 VSS.n2525 65.8183
R4804 VSS.t34 VSS.n2526 65.8183
R4805 VSS.t34 VSS.n2527 65.8183
R4806 VSS.t34 VSS.n2528 65.8183
R4807 VSS.t34 VSS.n2579 65.8183
R4808 VSS.t34 VSS.n2580 65.8183
R4809 VSS.t34 VSS.n2581 65.8183
R4810 VSS.t34 VSS.n2582 65.8183
R4811 VSS.t34 VSS.n2523 65.8183
R4812 VSS.t34 VSS.n2530 65.8183
R4813 VSS.t34 VSS.n2522 65.8183
R4814 VSS.t34 VSS.n2578 65.8183
R4815 VSS.t64 VSS.n2471 65.8183
R4816 VSS.t64 VSS.n2478 65.8183
R4817 VSS.t64 VSS.n2470 65.8183
R4818 VSS.t64 VSS.n2481 65.8183
R4819 VSS.t61 VSS.n2402 65.8183
R4820 VSS.t61 VSS.n2410 65.8183
R4821 VSS.t61 VSS.n2401 65.8183
R4822 VSS.t61 VSS.n2413 65.8183
R4823 VSS.t44 VSS.n1764 65.8183
R4824 VSS.t44 VSS.n1772 65.8183
R4825 VSS.t44 VSS.n1763 65.8183
R4826 VSS.n4630 VSS.t44 65.8183
R4827 VSS.t58 VSS.n1649 65.8183
R4828 VSS.t58 VSS.n1657 65.8183
R4829 VSS.t58 VSS.n1648 65.8183
R4830 VSS.t58 VSS.n1660 65.8183
R4831 VSS.t54 VSS.n2092 65.8183
R4832 VSS.t54 VSS.n2090 65.8183
R4833 VSS.t54 VSS.n2088 65.8183
R4834 VSS.t54 VSS.n2086 65.8183
R4835 VSS.n3270 VSS.t49 65.8183
R4836 VSS.n3238 VSS.t49 65.8183
R4837 VSS.n3240 VSS.t49 65.8183
R4838 VSS.n3366 VSS.t49 65.8183
R4839 VSS.t47 VSS.n2379 65.8183
R4840 VSS.t47 VSS.n2339 65.8183
R4841 VSS.t47 VSS.n2337 65.8183
R4842 VSS.t47 VSS.n2335 65.8183
R4843 VSS.n4394 VSS.t33 65.8183
R4844 VSS.n4397 VSS.t33 65.8183
R4845 VSS.n4399 VSS.t33 65.8183
R4846 VSS.n4619 VSS.t33 65.8183
R4847 VSS.t48 VSS.n1626 65.8183
R4848 VSS.t48 VSS.n1634 65.8183
R4849 VSS.t48 VSS.n1625 65.8183
R4850 VSS.t34 VSS.n2529 65.8183
R4851 VSS.t34 VSS.n2531 65.8183
R4852 VSS.t34 VSS.n2577 65.8183
R4853 VSS.t64 VSS.n2477 65.8183
R4854 VSS.t64 VSS.n2479 65.8183
R4855 VSS.t64 VSS.n2480 65.8183
R4856 VSS.t61 VSS.n2409 65.8183
R4857 VSS.t61 VSS.n2411 65.8183
R4858 VSS.t61 VSS.n2412 65.8183
R4859 VSS.t44 VSS.n1771 65.8183
R4860 VSS.t44 VSS.n1773 65.8183
R4861 VSS.t44 VSS.n1774 65.8183
R4862 VSS.t58 VSS.n1656 65.8183
R4863 VSS.t58 VSS.n1658 65.8183
R4864 VSS.t58 VSS.n1659 65.8183
R4865 VSS.t48 VSS.n1638 65.8183
R4866 VSS.t48 VSS.n1639 65.8183
R4867 VSS.t48 VSS.n1640 65.8183
R4868 VSS.t48 VSS.n1641 65.8183
R4869 VSS.t55 VSS.n1273 65.8183
R4870 VSS.t55 VSS.n1272 65.8183
R4871 VSS.t55 VSS.n1271 65.8183
R4872 VSS.t55 VSS.n1270 65.8183
R4873 VSS.t55 VSS.n1262 65.8183
R4874 VSS.t55 VSS.n1268 65.8183
R4875 VSS.t55 VSS.n1259 65.8183
R4876 VSS.t55 VSS.n1269 65.8183
R4877 VSS.t48 VSS.n1633 65.8183
R4878 VSS.t48 VSS.n1635 65.8183
R4879 VSS.t48 VSS.n1636 65.8183
R4880 VSS.n4716 VSS.t48 65.8183
R4881 VSS.t55 VSS.n1267 65.8183
R4882 VSS.t55 VSS.n1266 65.8183
R4883 VSS.t55 VSS.n1265 65.8183
R4884 VSS.t55 VSS.n1264 65.8183
R4885 VSS.t60 VSS.n1291 65.8183
R4886 VSS.t60 VSS.n1290 65.8183
R4887 VSS.t60 VSS.n1289 65.8183
R4888 VSS.t60 VSS.n1288 65.8183
R4889 VSS.t36 VSS.n88 65.8183
R4890 VSS.t36 VSS.n87 65.8183
R4891 VSS.t36 VSS.n82 65.8183
R4892 VSS.t36 VSS.n81 65.8183
R4893 VSS.t63 VSS.n384 65.8183
R4894 VSS.t63 VSS.n382 65.8183
R4895 VSS.t63 VSS.n381 65.8183
R4896 VSS.t63 VSS.n380 65.8183
R4897 VSS.n3498 VSS.t59 65.8183
R4898 VSS.n3496 VSS.t59 65.8183
R4899 VSS.n3469 VSS.t59 65.8183
R4900 VSS.n3902 VSS.t59 65.8183
R4901 VSS.t46 VSS.n769 65.8183
R4902 VSS.t46 VSS.n767 65.8183
R4903 VSS.t46 VSS.n766 65.8183
R4904 VSS.t46 VSS.n765 65.8183
R4905 VSS.t60 VSS.n1293 65.8183
R4906 VSS.t60 VSS.n1294 65.8183
R4907 VSS.n4764 VSS.t60 65.8183
R4908 VSS.t60 VSS.n4763 65.8183
R4909 VSS.t31 VSS.n115 65.8183
R4910 VSS.t31 VSS.n117 65.8183
R4911 VSS.t31 VSS.n118 65.8183
R4912 VSS.t56 VSS.n411 65.8183
R4913 VSS.t56 VSS.n413 65.8183
R4914 VSS.t56 VSS.n414 65.8183
R4915 VSS.t65 VSS.n2234 65.8183
R4916 VSS.t65 VSS.n2236 65.8183
R4917 VSS.t65 VSS.n2237 65.8183
R4918 VSS.t43 VSS.n796 65.8183
R4919 VSS.t43 VSS.n798 65.8183
R4920 VSS.t43 VSS.n799 65.8183
R4921 VSS.t55 VSS.n1263 65.8183
R4922 VSS.t55 VSS.n1261 65.8183
R4923 VSS.t55 VSS.n1260 65.8183
R4924 VSS.t55 VSS.n1258 65.8183
R4925 VSS.n480 VSS.t40 65.8183
R4926 VSS.n5517 VSS.t40 65.8183
R4927 VSS.n5507 VSS.t40 65.8183
R4928 VSS.n5224 VSS.t50 65.8183
R4929 VSS.n5211 VSS.t50 65.8183
R4930 VSS.n5209 VSS.t50 65.8183
R4931 VSS.n5270 VSS.t57 65.8183
R4932 VSS.n5257 VSS.t57 65.8183
R4933 VSS.n5255 VSS.t57 65.8183
R4934 VSS.n5316 VSS.t51 65.8183
R4935 VSS.n5303 VSS.t51 65.8183
R4936 VSS.n5301 VSS.t51 65.8183
R4937 VSS.t53 VSS.n928 65.8183
R4938 VSS.t53 VSS.n930 65.8183
R4939 VSS.t53 VSS.n931 65.8183
R4940 VSS.t62 VSS.n51 64.1729
R4941 VSS.t36 VSS.n90 64.1729
R4942 VSS.t46 VSS.n771 64.1729
R4943 VSS.n3529 VSS.t59 64.1729
R4944 VSS.t63 VSS.n386 64.1729
R4945 VSS.n3230 VSS.t49 64.1729
R4946 VSS.t54 VSS.n2094 64.1729
R4947 VSS.n1866 VSS.t33 64.1729
R4948 VSS.n3434 VSS.t47 64.1729
R4949 VSS.n3145 VSS.t34 64.1729
R4950 VSS.n3377 VSS.t64 64.1729
R4951 VSS.t61 VSS.n2408 64.1729
R4952 VSS.t44 VSS.n1770 64.1729
R4953 VSS.t58 VSS.n1655 64.1729
R4954 VSS.t48 VSS.n1632 64.1729
R4955 VSS.t31 VSS.n114 64.1729
R4956 VSS.t56 VSS.n410 64.1729
R4957 VSS.t65 VSS.n2233 64.1729
R4958 VSS.t43 VSS.n795 64.1729
R4959 VSS.n500 VSS.t40 64.1729
R4960 VSS.n5227 VSS.t50 64.1729
R4961 VSS.n5273 VSS.t57 64.1729
R4962 VSS.n5319 VSS.t51 64.1729
R4963 VSS.t53 VSS.n927 64.1729
R4964 VSS.n1512 VSS.n1511 62.4163
R4965 VSS.n4654 VSS.n1708 62.4163
R4966 VSS.n4199 VSS.n4076 62.4163
R4967 VSS.n4064 VSS.n128 62.4163
R4968 VSS.n4039 VSS.n4037 62.4163
R4969 VSS.n2600 VSS.n2599 62.4163
R4970 VSS.n4135 VSS.n4092 62.4163
R4971 VSS.n966 VSS.n869 62.4163
R4972 VSS.n183 VSS.n163 62.4163
R4973 VSS.n575 VSS.n229 62.4163
R4974 VSS.n5344 VSS.n5343 62.4163
R4975 VSS.n697 VSS.n676 62.4163
R4976 VSS.n4968 VSS.n699 62.4163
R4977 VSS.n997 VSS.n996 62.4163
R4978 VSS.n160 VSS.n158 62.4163
R4979 VSS.n3167 VSS.n2207 62.4163
R4980 VSS.n3417 VSS.n2215 62.4163
R4981 VSS.n660 VSS.n658 62.4163
R4982 VSS.n5054 VSS.n190 62.4163
R4983 VSS.n866 VSS.n864 62.4163
R4984 VSS.n2965 VSS.n2964 62.4163
R4985 VSS.n672 VSS.n669 62.4163
R4986 VSS.n2463 VSS.n2461 62.4163
R4987 VSS.n3001 VSS.n2905 62.4163
R4988 VSS.n4521 VSS.n1962 62.4163
R4989 VSS.n4527 VSS.n4526 62.4163
R4990 VSS.n2498 VSS.n2496 62.4163
R4991 VSS.t9 VSS.t23 60.0762
R4992 VSS.t23 VSS.t68 60.0762
R4993 VSS.t62 VSS.n22 57.8461
R4994 VSS.t36 VSS.n64 57.8461
R4995 VSS.t41 VSS.n358 57.8461
R4996 VSS.t60 VSS.n1615 57.8461
R4997 VSS.t45 VSS.n4832 57.8461
R4998 VSS.n4935 VSS.t42 57.8461
R4999 VSS.t46 VSS.n749 57.8461
R5000 VSS.n3847 VSS.t52 57.8461
R5001 VSS.n3882 VSS.t59 57.8461
R5002 VSS.t63 VSS.n367 57.8461
R5003 VSS.n3346 VSS.t49 57.8461
R5004 VSS.t54 VSS.n2099 57.8461
R5005 VSS.n4599 VSS.t33 57.8461
R5006 VSS.t47 VSS.n2386 57.8461
R5007 VSS.t34 VSS.n3144 57.8461
R5008 VSS.t64 VSS.n3376 57.8461
R5009 VSS.t61 VSS.n2397 57.8461
R5010 VSS.t44 VSS.n4629 57.8461
R5011 VSS.t58 VSS.n4711 57.8461
R5012 VSS.t31 VSS.n103 57.8461
R5013 VSS.t56 VSS.n399 57.8461
R5014 VSS.t65 VSS.n3912 57.8461
R5015 VSS.t43 VSS.n784 57.8461
R5016 VSS.t55 VSS.n4774 57.8461
R5017 VSS.n5494 VSS.t40 57.8461
R5018 VSS.n5196 VSS.t50 57.8461
R5019 VSS.n5242 VSS.t57 57.8461
R5020 VSS.n5288 VSS.t51 57.8461
R5021 VSS.t53 VSS.n4821 57.8461
R5022 VSS.n1922 VSS.n1632 56.6572
R5023 VSS.n1709 VSS.n1632 56.6572
R5024 VSS.n1820 VSS.n1655 56.6572
R5025 VSS.n2036 VSS.n1655 56.6572
R5026 VSS.n4428 VSS.n1770 56.6572
R5027 VSS.n4436 VSS.n1770 56.6572
R5028 VSS.n2896 VSS.n2408 56.6572
R5029 VSS.n2834 VSS.n2408 56.6572
R5030 VSS.n3378 VSS.n3377 56.6572
R5031 VSS.n3377 VSS.n2468 56.6572
R5032 VSS.n3501 VSS.n2233 56.6572
R5033 VSS.n3435 VSS.n3434 56.6572
R5034 VSS.n3434 VSS.n2334 56.6572
R5035 VSS.n3463 VSS.n2233 56.6572
R5036 VSS.n542 VSS.n90 56.6572
R5037 VSS.n455 VSS.n90 56.6572
R5038 VSS.n500 VSS.n499 56.6572
R5039 VSS.n458 VSS.n51 56.6572
R5040 VSS.n526 VSS.n51 56.6572
R5041 VSS.n501 VSS.n500 56.6572
R5042 VSS.n5227 VSS.n5226 56.6572
R5043 VSS.n5228 VSS.n5227 56.6572
R5044 VSS.n3750 VSS.n386 56.6572
R5045 VSS.n3748 VSS.n386 56.6572
R5046 VSS.n4795 VSS.n927 56.6572
R5047 VSS.n1324 VSS.n927 56.6572
R5048 VSS.n5319 VSS.n5318 56.6572
R5049 VSS.n5320 VSS.n5319 56.6572
R5050 VSS.n1122 VSS.n771 56.6572
R5051 VSS.n1120 VSS.n771 56.6572
R5052 VSS.n5273 VSS.n5272 56.6572
R5053 VSS.n5274 VSS.n5273 56.6572
R5054 VSS.n3530 VSS.n3529 56.6572
R5055 VSS.n3529 VSS.n3528 56.6572
R5056 VSS.n5386 VSS.n114 56.6572
R5057 VSS.n2148 VSS.n2094 56.6572
R5058 VSS.n2499 VSS.n2094 56.6572
R5059 VSS.n2152 VSS.n114 56.6572
R5060 VSS.n5093 VSS.n410 56.6572
R5061 VSS.n3315 VSS.n3230 56.6572
R5062 VSS.n3288 VSS.n3230 56.6572
R5063 VSS.n3291 VSS.n410 56.6572
R5064 VSS.n4865 VSS.n795 56.6572
R5065 VSS.n4568 VSS.n1866 56.6572
R5066 VSS.n4378 VSS.n1866 56.6572
R5067 VSS.n1869 VSS.n795 56.6572
R5068 VSS.n3146 VSS.n3145 56.6572
R5069 VSS.n3145 VSS.n2520 56.6572
R5070 VSS.n1244 VSS.n1219 56.3995
R5071 VSS.n1507 VSS.n1233 56.3995
R5072 VSS.n1511 VSS.n1233 56.3995
R5073 VSS.n1244 VSS.n1218 56.3995
R5074 VSS.n4134 VSS.n4090 56.3995
R5075 VSS.n4198 VSS.n4074 56.3995
R5076 VSS.n4225 VSS.n4224 56.3995
R5077 VSS.n4108 VSS.n12 56.3995
R5078 VSS.n2603 VSS.n2080 56.3995
R5079 VSS.n1731 VSS.n1728 56.3995
R5080 VSS.n2600 VSS.n2080 56.3995
R5081 VSS.n4224 VSS.n128 56.3995
R5082 VSS.n4199 VSS.n4198 56.3995
R5083 VSS.n4135 VSS.n4134 56.3995
R5084 VSS.n4109 VSS.n4108 56.3995
R5085 VSS.n1728 VSS.n1708 56.3995
R5086 VSS.n1486 VSS.n1485 56.3995
R5087 VSS.n4267 VSS.n4266 55.7181
R5088 VSS.n4281 VSS.n4267 55.7181
R5089 VSS.n4784 VSS.t32 55.7059
R5090 VSS.t32 VSS.n71 55.4806
R5091 VSS.t32 VSS.n29 55.4806
R5092 VSS.n1826 VSS.t32 55.4806
R5093 VSS.t45 VSS.n900 55.2026
R5094 VSS.t42 VSS.n737 55.2026
R5095 VSS.n3558 VSS.t52 55.2026
R5096 VSS.t41 VSS.n353 55.2026
R5097 VSS.n4775 VSS.t55 55.2026
R5098 VSS.t60 VSS.n1292 55.2026
R5099 VSS.n4283 VSS.n4282 54.5887
R5100 VSS.n4283 VSS.n4251 54.5887
R5101 VSS.t48 VSS.n1637 54.4705
R5102 VSS.n4720 VSS.n1269 53.3664
R5103 VSS.n1897 VSS.n1259 53.3664
R5104 VSS.n1938 VSS.n1268 53.3664
R5105 VSS.n1908 VSS.n1262 53.3664
R5106 VSS.n1451 VSS.n1264 53.3664
R5107 VSS.n1455 VSS.n1265 53.3664
R5108 VSS.n1459 VSS.n1266 53.3664
R5109 VSS.n1463 VSS.n1267 53.3664
R5110 VSS.n1275 VSS.n1258 53.3664
R5111 VSS.n1420 VSS.n1260 53.3664
R5112 VSS.n1435 VSS.n1261 53.3664
R5113 VSS.n1443 VSS.n1263 53.3664
R5114 VSS.n4724 VSS.n1273 53.3664
R5115 VSS.n4725 VSS.n1272 53.3664
R5116 VSS.n4729 VSS.n1271 53.3664
R5117 VSS.n4733 VSS.n1270 53.3664
R5118 VSS.n1643 VSS.n1625 53.3664
R5119 VSS.n1793 VSS.n1634 53.3664
R5120 VSS.n1804 VSS.n1626 53.3664
R5121 VSS.n4705 VSS.n1638 53.3664
R5122 VSS.n4701 VSS.n1639 53.3664
R5123 VSS.n4697 VSS.n1640 53.3664
R5124 VSS.n4693 VSS.n1641 53.3664
R5125 VSS.n4717 VSS.n4716 53.3664
R5126 VSS.n1899 VSS.n1636 53.3664
R5127 VSS.n1935 VSS.n1635 53.3664
R5128 VSS.n1913 VSS.n1633 53.3664
R5129 VSS.n1722 VSS.n1631 53.3664
R5130 VSS.n1718 VSS.n1630 53.3664
R5131 VSS.n1714 VSS.n1629 53.3664
R5132 VSS.n1710 VSS.n1628 53.3664
R5133 VSS.n1713 VSS.n1628 53.3664
R5134 VSS.n1717 VSS.n1629 53.3664
R5135 VSS.n1721 VSS.n1630 53.3664
R5136 VSS.n1724 VSS.n1631 53.3664
R5137 VSS.n2020 VSS.n1660 53.3664
R5138 VSS.n4357 VSS.n1648 53.3664
R5139 VSS.n4352 VSS.n1657 53.3664
R5140 VSS.n2033 VSS.n1649 53.3664
R5141 VSS.n2049 VSS.n1654 53.3664
R5142 VSS.n2045 VSS.n1653 53.3664
R5143 VSS.n2041 VSS.n1652 53.3664
R5144 VSS.n2037 VSS.n1651 53.3664
R5145 VSS.n2040 VSS.n1651 53.3664
R5146 VSS.n2044 VSS.n1652 53.3664
R5147 VSS.n2048 VSS.n1653 53.3664
R5148 VSS.n2051 VSS.n1654 53.3664
R5149 VSS.n1659 VSS.n1647 53.3664
R5150 VSS.n1800 VSS.n1658 53.3664
R5151 VSS.n1811 VSS.n1656 53.3664
R5152 VSS.n2016 VSS.n1661 53.3664
R5153 VSS.n2015 VSS.n1662 53.3664
R5154 VSS.n2011 VSS.n1663 53.3664
R5155 VSS.n2007 VSS.n1664 53.3664
R5156 VSS.n2019 VSS.n1661 53.3664
R5157 VSS.n2012 VSS.n1662 53.3664
R5158 VSS.n2008 VSS.n1663 53.3664
R5159 VSS.n1665 VSS.n1664 53.3664
R5160 VSS.n4631 VSS.n4630 53.3664
R5161 VSS.n4459 VSS.n1763 53.3664
R5162 VSS.n4474 VSS.n1772 53.3664
R5163 VSS.n4480 VSS.n1764 53.3664
R5164 VSS.n4449 VSS.n1769 53.3664
R5165 VSS.n4445 VSS.n1768 53.3664
R5166 VSS.n4441 VSS.n1767 53.3664
R5167 VSS.n4437 VSS.n1766 53.3664
R5168 VSS.n4440 VSS.n1766 53.3664
R5169 VSS.n4444 VSS.n1767 53.3664
R5170 VSS.n4448 VSS.n1768 53.3664
R5171 VSS.n4451 VSS.n1769 53.3664
R5172 VSS.n1828 VSS.n1774 53.3664
R5173 VSS.n4410 VSS.n1773 53.3664
R5174 VSS.n4419 VSS.n1771 53.3664
R5175 VSS.n2909 VSS.n1775 53.3664
R5176 VSS.n2910 VSS.n1776 53.3664
R5177 VSS.n2914 VSS.n1777 53.3664
R5178 VSS.n2918 VSS.n1778 53.3664
R5179 VSS.n1775 VSS.n1760 53.3664
R5180 VSS.n2913 VSS.n1776 53.3664
R5181 VSS.n2917 VSS.n1777 53.3664
R5182 VSS.n2920 VSS.n1778 53.3664
R5183 VSS.n2794 VSS.n2413 53.3664
R5184 VSS.n3049 VSS.n2401 53.3664
R5185 VSS.n3044 VSS.n2410 53.3664
R5186 VSS.n2807 VSS.n2402 53.3664
R5187 VSS.n2821 VSS.n2407 53.3664
R5188 VSS.n2825 VSS.n2406 53.3664
R5189 VSS.n2829 VSS.n2405 53.3664
R5190 VSS.n2833 VSS.n2404 53.3664
R5191 VSS.n2830 VSS.n2404 53.3664
R5192 VSS.n2826 VSS.n2405 53.3664
R5193 VSS.n2822 VSS.n2406 53.3664
R5194 VSS.n2818 VSS.n2407 53.3664
R5195 VSS.n2412 VSS.n2398 53.3664
R5196 VSS.n2878 VSS.n2411 53.3664
R5197 VSS.n2887 VSS.n2409 53.3664
R5198 VSS.n2790 VSS.n2414 53.3664
R5199 VSS.n2789 VSS.n2415 53.3664
R5200 VSS.n2785 VSS.n2416 53.3664
R5201 VSS.n3428 VSS.n3427 53.3664
R5202 VSS.n2793 VSS.n2414 53.3664
R5203 VSS.n2786 VSS.n2415 53.3664
R5204 VSS.n2418 VSS.n2416 53.3664
R5205 VSS.n3428 VSS.n2417 53.3664
R5206 VSS.n3090 VSS.n2481 53.3664
R5207 VSS.n2719 VSS.n2470 53.3664
R5208 VSS.n3079 VSS.n2478 53.3664
R5209 VSS.n2728 VSS.n2471 53.3664
R5210 VSS.n2742 VSS.n2476 53.3664
R5211 VSS.n2738 VSS.n2475 53.3664
R5212 VSS.n2734 VSS.n2474 53.3664
R5213 VSS.n2730 VSS.n2473 53.3664
R5214 VSS.n2733 VSS.n2473 53.3664
R5215 VSS.n2737 VSS.n2474 53.3664
R5216 VSS.n2741 VSS.n2475 53.3664
R5217 VSS.n2744 VSS.n2476 53.3664
R5218 VSS.n2490 VSS.n2480 53.3664
R5219 VSS.n3251 VSS.n2479 53.3664
R5220 VSS.n3260 VSS.n2477 53.3664
R5221 VSS.n2710 VSS.n2482 53.3664
R5222 VSS.n2709 VSS.n2483 53.3664
R5223 VSS.n2705 VSS.n2484 53.3664
R5224 VSS.n2701 VSS.n2485 53.3664
R5225 VSS.n3089 VSS.n2482 53.3664
R5226 VSS.n2706 VSS.n2483 53.3664
R5227 VSS.n2702 VSS.n2484 53.3664
R5228 VSS.n2698 VSS.n2485 53.3664
R5229 VSS.n3913 VSS.n2224 53.3664
R5230 VSS.n2226 VSS.n2222 53.3664
R5231 VSS.n2360 VSS.n2235 53.3664
R5232 VSS.n2367 VSS.n2227 53.3664
R5233 VSS.n2437 VSS.n2241 53.3664
R5234 VSS.n2436 VSS.n2240 53.3664
R5235 VSS.n2432 VSS.n2239 53.3664
R5236 VSS.n2428 VSS.n2238 53.3664
R5237 VSS.n2439 VSS.n2241 53.3664
R5238 VSS.n2433 VSS.n2240 53.3664
R5239 VSS.n2429 VSS.n2239 53.3664
R5240 VSS.n2425 VSS.n2238 53.3664
R5241 VSS.n2248 VSS.n2237 53.3664
R5242 VSS.n3481 VSS.n2236 53.3664
R5243 VSS.n3491 VSS.n2234 53.3664
R5244 VSS.n3450 VSS.n2232 53.3664
R5245 VSS.n3454 VSS.n2231 53.3664
R5246 VSS.n3458 VSS.n2230 53.3664
R5247 VSS.n3462 VSS.n2229 53.3664
R5248 VSS.n2392 VSS.n2335 53.3664
R5249 VSS.n2867 VSS.n2337 53.3664
R5250 VSS.n2859 VSS.n2339 53.3664
R5251 VSS.n2855 VSS.n2379 53.3664
R5252 VSS.n2456 VSS.n2387 53.3664
R5253 VSS.n2455 VSS.n2388 53.3664
R5254 VSS.n2451 VSS.n2389 53.3664
R5255 VSS.n2447 VSS.n2390 53.3664
R5256 VSS.n2391 VSS.n2387 53.3664
R5257 VSS.n2452 VSS.n2388 53.3664
R5258 VSS.n2448 VSS.n2389 53.3664
R5259 VSS.n2444 VSS.n2390 53.3664
R5260 VSS.n2384 VSS.n2336 53.3664
R5261 VSS.n2349 VSS.n2338 53.3664
R5262 VSS.n2378 VSS.n2340 53.3664
R5263 VSS.n2848 VSS.n2380 53.3664
R5264 VSS.n2844 VSS.n2381 53.3664
R5265 VSS.n2840 VSS.n2382 53.3664
R5266 VSS.n2836 VSS.n2383 53.3664
R5267 VSS.n2839 VSS.n2383 53.3664
R5268 VSS.n2843 VSS.n2382 53.3664
R5269 VSS.n2847 VSS.n2381 53.3664
R5270 VSS.n2851 VSS.n2380 53.3664
R5271 VSS.n3459 VSS.n2229 53.3664
R5272 VSS.n3455 VSS.n2230 53.3664
R5273 VSS.n3451 VSS.n2231 53.3664
R5274 VSS.n3447 VSS.n2232 53.3664
R5275 VSS.n100 VSS.n81 53.3664
R5276 VSS.n5403 VSS.n82 53.3664
R5277 VSS.n142 VSS.n87 53.3664
R5278 VSS.n5390 VSS.n88 53.3664
R5279 VSS.n4175 VSS.n95 53.3664
R5280 VSS.n4176 VSS.n96 53.3664
R5281 VSS.n4180 VSS.n97 53.3664
R5282 VSS.n4184 VSS.n98 53.3664
R5283 VSS.n99 VSS.n95 53.3664
R5284 VSS.n4179 VSS.n96 53.3664
R5285 VSS.n4183 VSS.n97 53.3664
R5286 VSS.n4187 VSS.n98 53.3664
R5287 VSS.n5452 VSS.n65 53.3664
R5288 VSS.n86 VSS.n85 53.3664
R5289 VSS.n5438 VSS.n5437 53.3664
R5290 VSS.n442 VSS.n91 53.3664
R5291 VSS.n446 VSS.n92 53.3664
R5292 VSS.n450 VSS.n93 53.3664
R5293 VSS.n454 VSS.n94 53.3664
R5294 VSS.n451 VSS.n94 53.3664
R5295 VSS.n447 VSS.n93 53.3664
R5296 VSS.n443 VSS.n92 53.3664
R5297 VSS.n439 VSS.n91 53.3664
R5298 VSS.n5477 VSS.n19 53.3664
R5299 VSS.n36 VSS.n35 53.3664
R5300 VSS.n5463 VSS.n5462 53.3664
R5301 VSS.n472 VSS.n38 53.3664
R5302 VSS.n5478 VSS.n17 53.3664
R5303 VSS.n5484 VSS.n5483 53.3664
R5304 VSS.n5487 VSS.n5486 53.3664
R5305 VSS.n5492 VSS.n5491 53.3664
R5306 VSS.n5479 VSS.n5478 53.3664
R5307 VSS.n5485 VSS.n5484 53.3664
R5308 VSS.n5486 VSS.n15 53.3664
R5309 VSS.n5493 VSS.n5492 53.3664
R5310 VSS.n5508 VSS.n5507 53.3664
R5311 VSS.n5517 VSS.n5516 53.3664
R5312 VSS.n480 VSS.n2 53.3664
R5313 VSS.n514 VSS.n513 53.3664
R5314 VSS.n509 VSS.n476 53.3664
R5315 VSS.n507 VSS.n506 53.3664
R5316 VSS.n502 VSS.n479 53.3664
R5317 VSS.n61 VSS.n42 53.3664
R5318 VSS.n74 VSS.n43 53.3664
R5319 VSS.n5441 VSS.n48 53.3664
R5320 VSS.n555 VSS.n49 53.3664
R5321 VSS.n4171 VSS.n56 53.3664
R5322 VSS.n4170 VSS.n57 53.3664
R5323 VSS.n4166 VSS.n58 53.3664
R5324 VSS.n4162 VSS.n59 53.3664
R5325 VSS.n60 VSS.n56 53.3664
R5326 VSS.n4167 VSS.n57 53.3664
R5327 VSS.n4163 VSS.n58 53.3664
R5328 VSS.n4159 VSS.n59 53.3664
R5329 VSS.n5473 VSS.n23 53.3664
R5330 VSS.n47 VSS.n46 53.3664
R5331 VSS.n5458 VSS.n5457 53.3664
R5332 VSS.n539 VSS.n52 53.3664
R5333 VSS.n535 VSS.n53 53.3664
R5334 VSS.n531 VSS.n54 53.3664
R5335 VSS.n527 VSS.n55 53.3664
R5336 VSS.n530 VSS.n55 53.3664
R5337 VSS.n534 VSS.n54 53.3664
R5338 VSS.n538 VSS.n53 53.3664
R5339 VSS.n558 VSS.n52 53.3664
R5340 VSS.n479 VSS.n477 53.3664
R5341 VSS.n508 VSS.n507 53.3664
R5342 VSS.n476 VSS.n474 53.3664
R5343 VSS.n515 VSS.n514 53.3664
R5344 VSS.n473 VSS.n472 53.3664
R5345 VSS.n5462 VSS.n5461 53.3664
R5346 VSS.n37 VSS.n36 53.3664
R5347 VSS.n34 VSS.n19 53.3664
R5348 VSS.n5457 VSS.n41 53.3664
R5349 VSS.n47 VSS.n40 53.3664
R5350 VSS.n45 VSS.n23 53.3664
R5351 VSS.n559 VSS.n49 53.3664
R5352 VSS.n554 VSS.n48 53.3664
R5353 VSS.n5442 VSS.n43 53.3664
R5354 VSS.n73 VSS.n42 53.3664
R5355 VSS.n5437 VSS.n80 53.3664
R5356 VSS.n86 VSS.n79 53.3664
R5357 VSS.n84 VSS.n65 53.3664
R5358 VSS.n5168 VSS.n335 53.3664
R5359 VSS.n5167 VSS.n341 53.3664
R5360 VSS.n3687 VSS.n3686 53.3664
R5361 VSS.n3709 VSS.n3708 53.3664
R5362 VSS.n3727 VSS.n3726 53.3664
R5363 VSS.n3722 VSS.n3714 53.3664
R5364 VSS.n3720 VSS.n3719 53.3664
R5365 VSS.n3715 VSS.n317 53.3664
R5366 VSS.n3716 VSS.n3715 53.3664
R5367 VSS.n3721 VSS.n3720 53.3664
R5368 VSS.n3714 VSS.n3712 53.3664
R5369 VSS.n3728 VSS.n3727 53.3664
R5370 VSS.n5209 VSS.n5208 53.3664
R5371 VSS.n5212 VSS.n5211 53.3664
R5372 VSS.n5224 VSS.n5223 53.3664
R5373 VSS.n5180 VSS.n5179 53.3664
R5374 VSS.n5182 VSS.n5181 53.3664
R5375 VSS.n5187 VSS.n5186 53.3664
R5376 VSS.n5190 VSS.n5189 53.3664
R5377 VSS.n5162 VSS.n5161 53.3664
R5378 VSS.n370 VSS.n356 53.3664
R5379 VSS.n5148 VSS.n355 53.3664
R5380 VSS.n3764 VSS.n354 53.3664
R5381 VSS.n3787 VSS.n349 53.3664
R5382 VSS.n3791 VSS.n350 53.3664
R5383 VSS.n3795 VSS.n351 53.3664
R5384 VSS.n3799 VSS.n352 53.3664
R5385 VSS.n5163 VSS.n345 53.3664
R5386 VSS.n346 VSS.n344 53.3664
R5387 VSS.n3691 VSS.n347 53.3664
R5388 VSS.n3704 VSS.n348 53.3664
R5389 VSS.n435 VSS.n359 53.3664
R5390 VSS.n434 VSS.n360 53.3664
R5391 VSS.n430 VSS.n361 53.3664
R5392 VSS.n426 VSS.n362 53.3664
R5393 VSS.n364 VSS.n359 53.3664
R5394 VSS.n431 VSS.n360 53.3664
R5395 VSS.n427 VSS.n361 53.3664
R5396 VSS.n423 VSS.n362 53.3664
R5397 VSS.n5179 VSS.n5178 53.3664
R5398 VSS.n5181 VSS.n333 53.3664
R5399 VSS.n5188 VSS.n5187 53.3664
R5400 VSS.n5189 VSS.n331 53.3664
R5401 VSS.n3710 VSS.n3709 53.3664
R5402 VSS.n3686 VSS.n3674 53.3664
R5403 VSS.n3685 VSS.n341 53.3664
R5404 VSS.n5169 VSS.n5168 53.3664
R5405 VSS.n3800 VSS.n348 53.3664
R5406 VSS.n3705 VSS.n347 53.3664
R5407 VSS.n3690 VSS.n346 53.3664
R5408 VSS.n5164 VSS.n5163 53.3664
R5409 VSS.n396 VSS.n380 53.3664
R5410 VSS.n5110 VSS.n381 53.3664
R5411 VSS.n642 VSS.n382 53.3664
R5412 VSS.n5097 VSS.n384 53.3664
R5413 VSS.n627 VSS.n391 53.3664
R5414 VSS.n626 VSS.n392 53.3664
R5415 VSS.n622 VSS.n393 53.3664
R5416 VSS.n618 VSS.n394 53.3664
R5417 VSS.n395 VSS.n391 53.3664
R5418 VSS.n623 VSS.n392 53.3664
R5419 VSS.n619 VSS.n393 53.3664
R5420 VSS.n615 VSS.n394 53.3664
R5421 VSS.n5157 VSS.n368 53.3664
R5422 VSS.n5144 VSS.n379 53.3664
R5423 VSS.n383 VSS.n377 53.3664
R5424 VSS.n3735 VSS.n387 53.3664
R5425 VSS.n3739 VSS.n388 53.3664
R5426 VSS.n3743 VSS.n389 53.3664
R5427 VSS.n3747 VSS.n390 53.3664
R5428 VSS.n3744 VSS.n390 53.3664
R5429 VSS.n3740 VSS.n389 53.3664
R5430 VSS.n3736 VSS.n388 53.3664
R5431 VSS.n3732 VSS.n387 53.3664
R5432 VSS.n3796 VSS.n352 53.3664
R5433 VSS.n3792 VSS.n351 53.3664
R5434 VSS.n3788 VSS.n350 53.3664
R5435 VSS.n3784 VSS.n349 53.3664
R5436 VSS.n1184 VSS.n932 53.3664
R5437 VSS.n4823 VSS.n4822 53.3664
R5438 VSS.n1351 VSS.n929 53.3664
R5439 VSS.n1348 VSS.n921 53.3664
R5440 VSS.n1188 VSS.n936 53.3664
R5441 VSS.n1189 VSS.n935 53.3664
R5442 VSS.n1193 VSS.n934 53.3664
R5443 VSS.n1197 VSS.n933 53.3664
R5444 VSS.n1185 VSS.n936 53.3664
R5445 VSS.n1192 VSS.n935 53.3664
R5446 VSS.n1196 VSS.n934 53.3664
R5447 VSS.n1199 VSS.n933 53.3664
R5448 VSS.n4812 VSS.n931 53.3664
R5449 VSS.n4808 VSS.n930 53.3664
R5450 VSS.n4800 VSS.n928 53.3664
R5451 VSS.n1337 VSS.n926 53.3664
R5452 VSS.n1333 VSS.n925 53.3664
R5453 VSS.n1329 VSS.n924 53.3664
R5454 VSS.n1325 VSS.n923 53.3664
R5455 VSS.n4834 VSS.n4833 53.3664
R5456 VSS.n1296 VSS.n895 53.3664
R5457 VSS.n1603 VSS.n905 53.3664
R5458 VSS.n1309 VSS.n898 53.3664
R5459 VSS.n1575 VSS.n901 53.3664
R5460 VSS.n1571 VSS.n902 53.3664
R5461 VSS.n1567 VSS.n903 53.3664
R5462 VSS.n1563 VSS.n904 53.3664
R5463 VSS.n911 VSS.n894 53.3664
R5464 VSS.n1358 VSS.n896 53.3664
R5465 VSS.n1367 VSS.n897 53.3664
R5466 VSS.n1376 VSS.n899 53.3664
R5467 VSS.n940 VSS.n909 53.3664
R5468 VSS.n941 VSS.n908 53.3664
R5469 VSS.n945 VSS.n907 53.3664
R5470 VSS.n949 VSS.n906 53.3664
R5471 VSS.n4763 VSS.n4762 53.3664
R5472 VSS.n4765 VSS.n4764 53.3664
R5473 VSS.n1413 VSS.n1294 53.3664
R5474 VSS.n1439 VSS.n1293 53.3664
R5475 VSS.n1474 VSS.n1288 53.3664
R5476 VSS.n1470 VSS.n1289 53.3664
R5477 VSS.n1466 VSS.n1290 53.3664
R5478 VSS.n1583 VSS.n1291 53.3664
R5479 VSS.n1613 VSS.n1284 53.3664
R5480 VSS.n1305 VSS.n1285 53.3664
R5481 VSS.n1598 VSS.n1286 53.3664
R5482 VSS.n1318 VSS.n1287 53.3664
R5483 VSS.n4758 VSS.n1616 53.3664
R5484 VSS.n4757 VSS.n1617 53.3664
R5485 VSS.n4753 VSS.n1618 53.3664
R5486 VSS.n4749 VSS.n1619 53.3664
R5487 VSS.n4761 VSS.n1616 53.3664
R5488 VSS.n4754 VSS.n1617 53.3664
R5489 VSS.n4750 VSS.n1618 53.3664
R5490 VSS.n4746 VSS.n1619 53.3664
R5491 VSS.n909 VSS.n892 53.3664
R5492 VSS.n944 VSS.n908 53.3664
R5493 VSS.n948 VSS.n907 53.3664
R5494 VSS.n951 VSS.n906 53.3664
R5495 VSS.n1587 VSS.n898 53.3664
R5496 VSS.n1308 VSS.n905 53.3664
R5497 VSS.n1602 VSS.n895 53.3664
R5498 VSS.n4833 VSS.n893 53.3664
R5499 VSS.n1584 VSS.n1287 53.3664
R5500 VSS.n1317 VSS.n1286 53.3664
R5501 VSS.n1599 VSS.n1285 53.3664
R5502 VSS.n1304 VSS.n1284 53.3664
R5503 VSS.n1566 VSS.n904 53.3664
R5504 VSS.n1570 VSS.n903 53.3664
R5505 VSS.n1574 VSS.n902 53.3664
R5506 VSS.n1578 VSS.n901 53.3664
R5507 VSS.n1328 VSS.n923 53.3664
R5508 VSS.n1332 VSS.n924 53.3664
R5509 VSS.n1336 VSS.n925 53.3664
R5510 VSS.n1339 VSS.n926 53.3664
R5511 VSS.n1344 VSS.n921 53.3664
R5512 VSS.n1349 VSS.n929 53.3664
R5513 VSS.n4822 VSS.n919 53.3664
R5514 VSS.n932 VSS.n918 53.3664
R5515 VSS.n1562 VSS.n899 53.3664
R5516 VSS.n1375 VSS.n897 53.3664
R5517 VSS.n1366 VSS.n896 53.3664
R5518 VSS.n1357 VSS.n894 53.3664
R5519 VSS.n4959 VSS.n4958 53.3664
R5520 VSS.n1043 VSS.n724 53.3664
R5521 VSS.n1070 VSS.n1069 53.3664
R5522 VSS.n1073 VSS.n1072 53.3664
R5523 VSS.n1100 VSS.n1099 53.3664
R5524 VSS.n1097 VSS.n1096 53.3664
R5525 VSS.n1092 VSS.n1089 53.3664
R5526 VSS.n1090 VSS.n279 53.3664
R5527 VSS.n1091 VSS.n1090 53.3664
R5528 VSS.n1089 VSS.n1087 53.3664
R5529 VSS.n1098 VSS.n1097 53.3664
R5530 VSS.n1101 VSS.n1100 53.3664
R5531 VSS.n5301 VSS.n5300 53.3664
R5532 VSS.n5304 VSS.n5303 53.3664
R5533 VSS.n5316 VSS.n5315 53.3664
R5534 VSS.n4955 VSS.n4954 53.3664
R5535 VSS.n4949 VSS.n4940 53.3664
R5536 VSS.n4948 VSS.n4947 53.3664
R5537 VSS.n4943 VSS.n4942 53.3664
R5538 VSS.n4934 VSS.n4933 53.3664
R5539 VSS.n752 VSS.n740 53.3664
R5540 VSS.n4920 VSS.n739 53.3664
R5541 VSS.n1136 VSS.n738 53.3664
R5542 VSS.n1159 VSS.n733 53.3664
R5543 VSS.n1163 VSS.n734 53.3664
R5544 VSS.n1167 VSS.n735 53.3664
R5545 VSS.n1171 VSS.n736 53.3664
R5546 VSS.n729 VSS.n728 53.3664
R5547 VSS.n1052 VSS.n730 53.3664
R5548 VSS.n1065 VSS.n731 53.3664
R5549 VSS.n1075 VSS.n732 53.3664
R5550 VSS.n817 VSS.n741 53.3664
R5551 VSS.n816 VSS.n742 53.3664
R5552 VSS.n812 VSS.n743 53.3664
R5553 VSS.n808 VSS.n744 53.3664
R5554 VSS.n746 VSS.n741 53.3664
R5555 VSS.n813 VSS.n742 53.3664
R5556 VSS.n809 VSS.n743 53.3664
R5557 VSS.n744 VSS.n726 53.3664
R5558 VSS.n4956 VSS.n4955 53.3664
R5559 VSS.n4950 VSS.n4949 53.3664
R5560 VSS.n4947 VSS.n4946 53.3664
R5561 VSS.n4942 VSS.n291 53.3664
R5562 VSS.n1072 VSS.n1038 53.3664
R5563 VSS.n1071 VSS.n1070 53.3664
R5564 VSS.n1044 VSS.n1043 53.3664
R5565 VSS.n4960 VSS.n4959 53.3664
R5566 VSS.n1170 VSS.n732 53.3664
R5567 VSS.n1076 VSS.n731 53.3664
R5568 VSS.n1066 VSS.n730 53.3664
R5569 VSS.n1051 VSS.n729 53.3664
R5570 VSS.n781 VSS.n765 53.3664
R5571 VSS.n4882 VSS.n766 53.3664
R5572 VSS.n849 VSS.n767 53.3664
R5573 VSS.n4869 VSS.n769 53.3664
R5574 VSS.n835 VSS.n776 53.3664
R5575 VSS.n834 VSS.n777 53.3664
R5576 VSS.n830 VSS.n778 53.3664
R5577 VSS.n826 VSS.n779 53.3664
R5578 VSS.n780 VSS.n776 53.3664
R5579 VSS.n831 VSS.n777 53.3664
R5580 VSS.n827 VSS.n778 53.3664
R5581 VSS.n823 VSS.n779 53.3664
R5582 VSS.n4929 VSS.n750 53.3664
R5583 VSS.n4916 VSS.n764 53.3664
R5584 VSS.n768 VSS.n762 53.3664
R5585 VSS.n1107 VSS.n772 53.3664
R5586 VSS.n1111 VSS.n773 53.3664
R5587 VSS.n1115 VSS.n774 53.3664
R5588 VSS.n1119 VSS.n775 53.3664
R5589 VSS.n1116 VSS.n775 53.3664
R5590 VSS.n1112 VSS.n774 53.3664
R5591 VSS.n1108 VSS.n773 53.3664
R5592 VSS.n1104 VSS.n772 53.3664
R5593 VSS.n1168 VSS.n736 53.3664
R5594 VSS.n1164 VSS.n735 53.3664
R5595 VSS.n1160 VSS.n734 53.3664
R5596 VSS.n1156 VSS.n733 53.3664
R5597 VSS.n1144 VSS.n738 53.3664
R5598 VSS.n1135 VSS.n739 53.3664
R5599 VSS.n4921 VSS.n740 53.3664
R5600 VSS.n4934 VSS.n745 53.3664
R5601 VSS.n1126 VSS.n768 53.3664
R5602 VSS.n4917 VSS.n4916 53.3664
R5603 VSS.n763 VSS.n750 53.3664
R5604 VSS.n3831 VSS.n3830 53.3664
R5605 VSS.n3835 VSS.n3834 53.3664
R5606 VSS.n3629 VSS.n2283 53.3664
R5607 VSS.n3612 VSS.n3611 53.3664
R5608 VSS.n3597 VSS.n3584 53.3664
R5609 VSS.n3595 VSS.n3594 53.3664
R5610 VSS.n3590 VSS.n3587 53.3664
R5611 VSS.n3588 VSS.n298 53.3664
R5612 VSS.n3589 VSS.n3588 53.3664
R5613 VSS.n3587 VSS.n3585 53.3664
R5614 VSS.n3596 VSS.n3595 53.3664
R5615 VSS.n3584 VSS.n2296 53.3664
R5616 VSS.n5255 VSS.n5254 53.3664
R5617 VSS.n5258 VSS.n5257 53.3664
R5618 VSS.n5270 VSS.n5269 53.3664
R5619 VSS.n3828 VSS.n3827 53.3664
R5620 VSS.n3822 VSS.n3813 53.3664
R5621 VSS.n3821 VSS.n3820 53.3664
R5622 VSS.n3816 VSS.n3815 53.3664
R5623 VSS.n3866 VSS.n3865 53.3664
R5624 VSS.n3870 VSS.n3869 53.3664
R5625 VSS.n2313 VSS.n2265 53.3664
R5626 VSS.n3556 VSS.n3555 53.3664
R5627 VSS.n3572 VSS.n3571 53.3664
R5628 VSS.n3573 VSS.n2305 53.3664
R5629 VSS.n3580 VSS.n3579 53.3664
R5630 VSS.n3602 VSS.n2303 53.3664
R5631 VSS.n3622 VSS.n2274 53.3664
R5632 VSS.n3625 VSS.n3624 53.3664
R5633 VSS.n3621 VSS.n2285 53.3664
R5634 VSS.n3605 VSS.n3604 53.3664
R5635 VSS.n3863 VSS.n3862 53.3664
R5636 VSS.n3857 VSS.n2270 53.3664
R5637 VSS.n3856 VSS.n3855 53.3664
R5638 VSS.n3849 VSS.n2272 53.3664
R5639 VSS.n3864 VSS.n3863 53.3664
R5640 VSS.n3858 VSS.n3857 53.3664
R5641 VSS.n3855 VSS.n3854 53.3664
R5642 VSS.n3850 VSS.n3849 53.3664
R5643 VSS.n3829 VSS.n3828 53.3664
R5644 VSS.n3823 VSS.n3822 53.3664
R5645 VSS.n3820 VSS.n3819 53.3664
R5646 VSS.n3815 VSS.n310 53.3664
R5647 VSS.n3613 VSS.n3612 53.3664
R5648 VSS.n3610 VSS.n2283 53.3664
R5649 VSS.n3836 VSS.n3835 53.3664
R5650 VSS.n3832 VSS.n3831 53.3664
R5651 VSS.n3606 VSS.n3605 53.3664
R5652 VSS.n3603 VSS.n2285 53.3664
R5653 VSS.n3626 VSS.n3625 53.3664
R5654 VSS.n3623 VSS.n3622 53.3664
R5655 VSS.n3902 VSS.n3901 53.3664
R5656 VSS.n3469 VSS.n2250 53.3664
R5657 VSS.n3496 VSS.n3495 53.3664
R5658 VSS.n3499 VSS.n3498 53.3664
R5659 VSS.n3898 VSS.n3897 53.3664
R5660 VSS.n3892 VSS.n2252 53.3664
R5661 VSS.n3891 VSS.n3890 53.3664
R5662 VSS.n3884 VSS.n2254 53.3664
R5663 VSS.n3899 VSS.n3898 53.3664
R5664 VSS.n3893 VSS.n3892 53.3664
R5665 VSS.n3890 VSS.n3889 53.3664
R5666 VSS.n3885 VSS.n3884 53.3664
R5667 VSS.n3532 VSS.n2256 53.3664
R5668 VSS.n3535 VSS.n3534 53.3664
R5669 VSS.n3551 VSS.n3550 53.3664
R5670 VSS.n3515 VSS.n3514 53.3664
R5671 VSS.n3516 VSS.n2319 53.3664
R5672 VSS.n3523 VSS.n3522 53.3664
R5673 VSS.n3527 VSS.n2317 53.3664
R5674 VSS.n3524 VSS.n2317 53.3664
R5675 VSS.n3522 VSS.n3521 53.3664
R5676 VSS.n3517 VSS.n3516 53.3664
R5677 VSS.n3514 VSS.n3513 53.3664
R5678 VSS.n3581 VSS.n2303 53.3664
R5679 VSS.n3579 VSS.n3578 53.3664
R5680 VSS.n3574 VSS.n3573 53.3664
R5681 VSS.n3571 VSS.n3570 53.3664
R5682 VSS.n3557 VSS.n3556 53.3664
R5683 VSS.n2314 VSS.n2313 53.3664
R5684 VSS.n3871 VSS.n3870 53.3664
R5685 VSS.n3867 VSS.n3866 53.3664
R5686 VSS.n3552 VSS.n3551 53.3664
R5687 VSS.n3536 VSS.n3535 53.3664
R5688 VSS.n3533 VSS.n3532 53.3664
R5689 VSS.n3772 VSS.n354 53.3664
R5690 VSS.n3763 VSS.n355 53.3664
R5691 VSS.n5149 VSS.n356 53.3664
R5692 VSS.n5162 VSS.n363 53.3664
R5693 VSS.n3754 VSS.n383 53.3664
R5694 VSS.n5145 VSS.n5144 53.3664
R5695 VSS.n378 VSS.n368 53.3664
R5696 VSS.n2116 VSS.n119 53.3664
R5697 VSS.n3990 VSS.n107 53.3664
R5698 VSS.n2128 VSS.n116 53.3664
R5699 VSS.n3977 VSS.n108 53.3664
R5700 VSS.n5431 VSS.n5430 53.3664
R5701 VSS.n124 VSS.n122 53.3664
R5702 VSS.n5425 VSS.n121 53.3664
R5703 VSS.n5421 VSS.n120 53.3664
R5704 VSS.n5431 VSS.n123 53.3664
R5705 VSS.n5426 VSS.n122 53.3664
R5706 VSS.n5422 VSS.n121 53.3664
R5707 VSS.n5418 VSS.n120 53.3664
R5708 VSS.n118 VSS.n104 53.3664
R5709 VSS.n5399 VSS.n117 53.3664
R5710 VSS.n146 VSS.n115 53.3664
R5711 VSS.n2165 VSS.n113 53.3664
R5712 VSS.n2161 VSS.n112 53.3664
R5713 VSS.n2157 VSS.n111 53.3664
R5714 VSS.n2153 VSS.n110 53.3664
R5715 VSS.n2086 VSS.n2085 53.3664
R5716 VSS.n2542 VSS.n2088 53.3664
R5717 VSS.n2567 VSS.n2090 53.3664
R5718 VSS.n2554 VSS.n2092 53.3664
R5719 VSS.n2106 VSS.n2100 53.3664
R5720 VSS.n2107 VSS.n2101 53.3664
R5721 VSS.n2111 VSS.n2102 53.3664
R5722 VSS.n4004 VSS.n4003 53.3664
R5723 VSS.n2100 VSS.n2084 53.3664
R5724 VSS.n2110 VSS.n2101 53.3664
R5725 VSS.n2104 VSS.n2102 53.3664
R5726 VSS.n4004 VSS.n2103 53.3664
R5727 VSS.n2122 VSS.n2087 53.3664
R5728 VSS.n3986 VSS.n2089 53.3664
R5729 VSS.n2137 VSS.n2091 53.3664
R5730 VSS.n2512 VSS.n2095 53.3664
R5731 VSS.n2508 VSS.n2096 53.3664
R5732 VSS.n2504 VSS.n2097 53.3664
R5733 VSS.n2500 VSS.n2098 53.3664
R5734 VSS.n2503 VSS.n2098 53.3664
R5735 VSS.n2507 VSS.n2097 53.3664
R5736 VSS.n2511 VSS.n2096 53.3664
R5737 VSS.n2516 VSS.n2095 53.3664
R5738 VSS.n2156 VSS.n110 53.3664
R5739 VSS.n2160 VSS.n111 53.3664
R5740 VSS.n2164 VSS.n112 53.3664
R5741 VSS.n2167 VSS.n113 53.3664
R5742 VSS.n3200 VSS.n415 53.3664
R5743 VSS.n3211 VSS.n403 53.3664
R5744 VSS.n3334 VSS.n412 53.3664
R5745 VSS.n3219 VSS.n404 53.3664
R5746 VSS.n5138 VSS.n5137 53.3664
R5747 VSS.n420 VSS.n418 53.3664
R5748 VSS.n5132 VSS.n417 53.3664
R5749 VSS.n5128 VSS.n416 53.3664
R5750 VSS.n5138 VSS.n419 53.3664
R5751 VSS.n5133 VSS.n418 53.3664
R5752 VSS.n5129 VSS.n417 53.3664
R5753 VSS.n5125 VSS.n416 53.3664
R5754 VSS.n414 VSS.n400 53.3664
R5755 VSS.n5106 VSS.n413 53.3664
R5756 VSS.n646 VSS.n411 53.3664
R5757 VSS.n3304 VSS.n409 53.3664
R5758 VSS.n3300 VSS.n408 53.3664
R5759 VSS.n3296 VSS.n407 53.3664
R5760 VSS.n3292 VSS.n406 53.3664
R5761 VSS.n3366 VSS.n3365 53.3664
R5762 VSS.n3240 VSS.n2492 53.3664
R5763 VSS.n3239 VSS.n3238 53.3664
R5764 VSS.n3270 VSS.n3269 53.3664
R5765 VSS.n3362 VSS.n3361 53.3664
R5766 VSS.n3356 VSS.n3195 53.3664
R5767 VSS.n3355 VSS.n3354 53.3664
R5768 VSS.n3348 VSS.n3197 53.3664
R5769 VSS.n3363 VSS.n3362 53.3664
R5770 VSS.n3357 VSS.n3356 53.3664
R5771 VSS.n3354 VSS.n3353 53.3664
R5772 VSS.n3349 VSS.n3348 53.3664
R5773 VSS.n3327 VSS.n3199 53.3664
R5774 VSS.n3330 VSS.n3329 53.3664
R5775 VSS.n3326 VSS.n3216 53.3664
R5776 VSS.n3274 VSS.n3273 53.3664
R5777 VSS.n3279 VSS.n3278 53.3664
R5778 VSS.n3280 VSS.n3233 53.3664
R5779 VSS.n3287 VSS.n3286 53.3664
R5780 VSS.n3286 VSS.n3285 53.3664
R5781 VSS.n3281 VSS.n3280 53.3664
R5782 VSS.n3278 VSS.n3277 53.3664
R5783 VSS.n3273 VSS.n3272 53.3664
R5784 VSS.n3295 VSS.n406 53.3664
R5785 VSS.n3299 VSS.n407 53.3664
R5786 VSS.n3303 VSS.n408 53.3664
R5787 VSS.n3306 VSS.n409 53.3664
R5788 VSS.n3318 VSS.n404 53.3664
R5789 VSS.n3218 VSS.n412 53.3664
R5790 VSS.n3335 VSS.n403 53.3664
R5791 VSS.n3210 VSS.n415 53.3664
R5792 VSS.n3229 VSS.n3216 53.3664
R5793 VSS.n3331 VSS.n3330 53.3664
R5794 VSS.n3328 VSS.n3327 53.3664
R5795 VSS.n2140 VSS.n108 53.3664
R5796 VSS.n3978 VSS.n116 53.3664
R5797 VSS.n2127 VSS.n107 53.3664
R5798 VSS.n3991 VSS.n119 53.3664
R5799 VSS.n3974 VSS.n2091 53.3664
R5800 VSS.n2136 VSS.n2089 53.3664
R5801 VSS.n3987 VSS.n2087 53.3664
R5802 VSS.n1837 VSS.n800 53.3664
R5803 VSS.n1847 VSS.n788 53.3664
R5804 VSS.n4587 VSS.n797 53.3664
R5805 VSS.n1855 VSS.n789 53.3664
R5806 VSS.n4910 VSS.n4909 53.3664
R5807 VSS.n805 VSS.n803 53.3664
R5808 VSS.n4904 VSS.n802 53.3664
R5809 VSS.n4900 VSS.n801 53.3664
R5810 VSS.n4910 VSS.n804 53.3664
R5811 VSS.n4905 VSS.n803 53.3664
R5812 VSS.n4901 VSS.n802 53.3664
R5813 VSS.n4897 VSS.n801 53.3664
R5814 VSS.n799 VSS.n785 53.3664
R5815 VSS.n4878 VSS.n798 53.3664
R5816 VSS.n853 VSS.n796 53.3664
R5817 VSS.n1882 VSS.n794 53.3664
R5818 VSS.n1878 VSS.n793 53.3664
R5819 VSS.n1874 VSS.n792 53.3664
R5820 VSS.n1870 VSS.n791 53.3664
R5821 VSS.n4619 VSS.n4618 53.3664
R5822 VSS.n4399 VSS.n1830 53.3664
R5823 VSS.n4398 VSS.n4397 53.3664
R5824 VSS.n4395 VSS.n4394 53.3664
R5825 VSS.n4615 VSS.n4614 53.3664
R5826 VSS.n4609 VSS.n1832 53.3664
R5827 VSS.n4608 VSS.n4607 53.3664
R5828 VSS.n4601 VSS.n1834 53.3664
R5829 VSS.n4616 VSS.n4615 53.3664
R5830 VSS.n4610 VSS.n4609 53.3664
R5831 VSS.n4607 VSS.n4606 53.3664
R5832 VSS.n4602 VSS.n4601 53.3664
R5833 VSS.n4580 VSS.n1836 53.3664
R5834 VSS.n4583 VSS.n4582 53.3664
R5835 VSS.n4579 VSS.n1852 53.3664
R5836 VSS.n4391 VSS.n4390 53.3664
R5837 VSS.n4386 VSS.n4374 53.3664
R5838 VSS.n4384 VSS.n4383 53.3664
R5839 VSS.n4379 VSS.n4377 53.3664
R5840 VSS.n4377 VSS.n4375 53.3664
R5841 VSS.n4385 VSS.n4384 53.3664
R5842 VSS.n4374 VSS.n4372 53.3664
R5843 VSS.n4392 VSS.n4391 53.3664
R5844 VSS.n1873 VSS.n791 53.3664
R5845 VSS.n1877 VSS.n792 53.3664
R5846 VSS.n1881 VSS.n793 53.3664
R5847 VSS.n1884 VSS.n794 53.3664
R5848 VSS.n4571 VSS.n789 53.3664
R5849 VSS.n1854 VSS.n797 53.3664
R5850 VSS.n4588 VSS.n788 53.3664
R5851 VSS.n1846 VSS.n800 53.3664
R5852 VSS.n1865 VSS.n1852 53.3664
R5853 VSS.n4584 VSS.n4583 53.3664
R5854 VSS.n4581 VSS.n4580 53.3664
R5855 VSS.n2342 VSS.n2227 53.3664
R5856 VSS.n2368 VSS.n2235 53.3664
R5857 VSS.n2359 VSS.n2226 53.3664
R5858 VSS.n3914 VSS.n3913 53.3664
R5859 VSS.n2378 VSS.n2377 53.3664
R5860 VSS.n2347 VSS.n2338 53.3664
R5861 VSS.n2350 VSS.n2336 53.3664
R5862 VSS.n3125 VSS.n2578 53.3664
R5863 VSS.n2632 VSS.n2522 53.3664
R5864 VSS.n3114 VSS.n2530 53.3664
R5865 VSS.n2641 VSS.n2523 53.3664
R5866 VSS.n2655 VSS.n2528 53.3664
R5867 VSS.n2651 VSS.n2527 53.3664
R5868 VSS.n2647 VSS.n2526 53.3664
R5869 VSS.n2643 VSS.n2525 53.3664
R5870 VSS.n2646 VSS.n2525 53.3664
R5871 VSS.n2650 VSS.n2526 53.3664
R5872 VSS.n2654 VSS.n2527 53.3664
R5873 VSS.n2657 VSS.n2528 53.3664
R5874 VSS.n2577 VSS.n2576 53.3664
R5875 VSS.n2545 VSS.n2531 53.3664
R5876 VSS.n2563 VSS.n2529 53.3664
R5877 VSS.n3129 VSS.n2579 53.3664
R5878 VSS.n3130 VSS.n2580 53.3664
R5879 VSS.n3134 VSS.n2581 53.3664
R5880 VSS.n3138 VSS.n2582 53.3664
R5881 VSS.n3126 VSS.n2579 53.3664
R5882 VSS.n3133 VSS.n2580 53.3664
R5883 VSS.n3137 VSS.n2581 53.3664
R5884 VSS.n3141 VSS.n2582 53.3664
R5885 VSS.n3104 VSS.n2523 53.3664
R5886 VSS.n2640 VSS.n2530 53.3664
R5887 VSS.n3115 VSS.n2522 53.3664
R5888 VSS.n2631 VSS.n2578 53.3664
R5889 VSS.n3069 VSS.n2471 53.3664
R5890 VSS.n2727 VSS.n2478 53.3664
R5891 VSS.n3080 VSS.n2470 53.3664
R5892 VSS.n2718 VSS.n2481 53.3664
R5893 VSS.n3034 VSS.n2402 53.3664
R5894 VSS.n2806 VSS.n2410 53.3664
R5895 VSS.n3045 VSS.n2401 53.3664
R5896 VSS.n3048 VSS.n2413 53.3664
R5897 VSS.n4453 VSS.n1764 53.3664
R5898 VSS.n4479 VSS.n1772 53.3664
R5899 VSS.n4473 VSS.n1763 53.3664
R5900 VSS.n4630 VSS.n1761 53.3664
R5901 VSS.n4342 VSS.n1649 53.3664
R5902 VSS.n2032 VSS.n1657 53.3664
R5903 VSS.n4353 VSS.n1648 53.3664
R5904 VSS.n4356 VSS.n1660 53.3664
R5905 VSS.n2517 VSS.n2092 53.3664
R5906 VSS.n2553 VSS.n2090 53.3664
R5907 VSS.n2568 VSS.n2088 53.3664
R5908 VSS.n2541 VSS.n2086 53.3664
R5909 VSS.n3271 VSS.n3270 53.3664
R5910 VSS.n3238 VSS.n3235 53.3664
R5911 VSS.n3241 VSS.n3240 53.3664
R5912 VSS.n3367 VSS.n3366 53.3664
R5913 VSS.n2852 VSS.n2379 53.3664
R5914 VSS.n2856 VSS.n2339 53.3664
R5915 VSS.n2860 VSS.n2337 53.3664
R5916 VSS.n2868 VSS.n2335 53.3664
R5917 VSS.n4394 VSS.n4393 53.3664
R5918 VSS.n4397 VSS.n4396 53.3664
R5919 VSS.n4400 VSS.n4399 53.3664
R5920 VSS.n4620 VSS.n4619 53.3664
R5921 VSS.n1814 VSS.n1626 53.3664
R5922 VSS.n1805 VSS.n1634 53.3664
R5923 VSS.n1794 VSS.n1625 53.3664
R5924 VSS.n2529 VSS.n2519 53.3664
R5925 VSS.n2564 VSS.n2531 53.3664
R5926 VSS.n2577 VSS.n2532 53.3664
R5927 VSS.n2477 VSS.n2467 53.3664
R5928 VSS.n3259 VSS.n2479 53.3664
R5929 VSS.n3250 VSS.n2480 53.3664
R5930 VSS.n2895 VSS.n2409 53.3664
R5931 VSS.n2886 VSS.n2411 53.3664
R5932 VSS.n2877 VSS.n2412 53.3664
R5933 VSS.n4427 VSS.n1771 53.3664
R5934 VSS.n4418 VSS.n1773 53.3664
R5935 VSS.n4409 VSS.n1774 53.3664
R5936 VSS.n1819 VSS.n1656 53.3664
R5937 VSS.n1810 VSS.n1658 53.3664
R5938 VSS.n1799 VSS.n1659 53.3664
R5939 VSS.n4702 VSS.n1638 53.3664
R5940 VSS.n4698 VSS.n1639 53.3664
R5941 VSS.n4694 VSS.n1640 53.3664
R5942 VSS.n1641 VSS.n1623 53.3664
R5943 VSS.n4721 VSS.n1273 53.3664
R5944 VSS.n4728 VSS.n1272 53.3664
R5945 VSS.n4732 VSS.n1271 53.3664
R5946 VSS.n4735 VSS.n1270 53.3664
R5947 VSS.n1925 VSS.n1262 53.3664
R5948 VSS.n1909 VSS.n1268 53.3664
R5949 VSS.n1939 VSS.n1259 53.3664
R5950 VSS.n1896 VSS.n1269 53.3664
R5951 VSS.n1923 VSS.n1633 53.3664
R5952 VSS.n1912 VSS.n1635 53.3664
R5953 VSS.n1934 VSS.n1636 53.3664
R5954 VSS.n4716 VSS.n1624 53.3664
R5955 VSS.n1460 VSS.n1267 53.3664
R5956 VSS.n1456 VSS.n1266 53.3664
R5957 VSS.n1452 VSS.n1265 53.3664
R5958 VSS.n1264 VSS.n1256 53.3664
R5959 VSS.n1465 VSS.n1291 53.3664
R5960 VSS.n1469 VSS.n1290 53.3664
R5961 VSS.n1473 VSS.n1289 53.3664
R5962 VSS.n1477 VSS.n1288 53.3664
R5963 VSS.n438 VSS.n88 53.3664
R5964 VSS.n5391 VSS.n87 53.3664
R5965 VSS.n141 VSS.n82 53.3664
R5966 VSS.n5404 VSS.n81 53.3664
R5967 VSS.n3731 VSS.n384 53.3664
R5968 VSS.n5098 VSS.n382 53.3664
R5969 VSS.n641 VSS.n381 53.3664
R5970 VSS.n5111 VSS.n380 53.3664
R5971 VSS.n3498 VSS.n2321 53.3664
R5972 VSS.n3497 VSS.n3496 53.3664
R5973 VSS.n3470 VSS.n3469 53.3664
R5974 VSS.n3903 VSS.n3902 53.3664
R5975 VSS.n1103 VSS.n769 53.3664
R5976 VSS.n4870 VSS.n767 53.3664
R5977 VSS.n848 VSS.n766 53.3664
R5978 VSS.n4883 VSS.n765 53.3664
R5979 VSS.n1446 VSS.n1293 53.3664
R5980 VSS.n1438 VSS.n1294 53.3664
R5981 VSS.n4764 VSS.n1283 53.3664
R5982 VSS.n4763 VSS.n1282 53.3664
R5983 VSS.n5387 VSS.n115 53.3664
R5984 VSS.n145 VSS.n117 53.3664
R5985 VSS.n5400 VSS.n118 53.3664
R5986 VSS.n5094 VSS.n411 53.3664
R5987 VSS.n645 VSS.n413 53.3664
R5988 VSS.n5107 VSS.n414 53.3664
R5989 VSS.n3502 VSS.n2234 53.3664
R5990 VSS.n3492 VSS.n2236 53.3664
R5991 VSS.n3480 VSS.n2237 53.3664
R5992 VSS.n4866 VSS.n796 53.3664
R5993 VSS.n852 VSS.n798 53.3664
R5994 VSS.n4879 VSS.n799 53.3664
R5995 VSS.n1462 VSS.n1263 53.3664
R5996 VSS.n1442 VSS.n1261 53.3664
R5997 VSS.n1434 VSS.n1260 53.3664
R5998 VSS.n1419 VSS.n1258 53.3664
R5999 VSS.n481 VSS.n480 53.3664
R6000 VSS.n5518 VSS.n5517 53.3664
R6001 VSS.n5507 VSS.n3 53.3664
R6002 VSS.n5225 VSS.n5224 53.3664
R6003 VSS.n5211 VSS.n320 53.3664
R6004 VSS.n5210 VSS.n5209 53.3664
R6005 VSS.n5271 VSS.n5270 53.3664
R6006 VSS.n5257 VSS.n301 53.3664
R6007 VSS.n5256 VSS.n5255 53.3664
R6008 VSS.n5317 VSS.n5316 53.3664
R6009 VSS.n5303 VSS.n282 53.3664
R6010 VSS.n5302 VSS.n5301 53.3664
R6011 VSS.n4796 VSS.n928 53.3664
R6012 VSS.n4799 VSS.n930 53.3664
R6013 VSS.n4809 VSS.n931 53.3664
R6014 VSS.n4268 VSS.t69 52.4309
R6015 VSS.n4252 VSS.t90 52.242
R6016 VSS.n183 VSS.n180 49.7381
R6017 VSS.n190 VSS.n184 49.7381
R6018 VSS.n697 VSS.n185 49.7381
R6019 VSS.n966 VSS.n186 49.7381
R6020 VSS.n229 VSS.n223 49.7381
R6021 VSS.n5343 VSS.n5342 49.7381
R6022 VSS.n4968 VSS.n224 49.7381
R6023 VSS.n997 VSS.n225 49.7381
R6024 VSS.n630 VSS.n160 49.7381
R6025 VSS.n5052 VSS.n660 49.7381
R6026 VSS.n669 VSS.n664 49.7381
R6027 VSS.n866 VSS.n665 49.7381
R6028 VSS.n2209 VSS.n2207 49.7381
R6029 VSS.n2215 VSS.n2210 49.7381
R6030 VSS.n2964 VSS.n2211 49.7381
R6031 VSS.n4527 VSS.n1952 49.7381
R6032 VSS.n2498 VSS.n2497 49.7381
R6033 VSS.n2463 VSS.n2462 49.7381
R6034 VSS.n2928 VSS.n2905 49.7381
R6035 VSS.n4522 VSS.n1962 49.7381
R6036 VSS.n5361 VSS.n183 48.7629
R6037 VSS.n5359 VSS.n190 48.7629
R6038 VSS.n697 VSS.n188 48.7629
R6039 VSS.n966 VSS.n187 48.7629
R6040 VSS.n5340 VSS.n229 48.7629
R6041 VSS.n5343 VSS.n221 48.7629
R6042 VSS.n4968 VSS.n227 48.7629
R6043 VSS.n997 VSS.n226 48.7629
R6044 VSS.n160 VSS.n156 48.7629
R6045 VSS.n660 VSS.n656 48.7629
R6046 VSS.n5050 VSS.n669 48.7629
R6047 VSS.n866 VSS.n667 48.7629
R6048 VSS.n3962 VSS.n2207 48.7629
R6049 VSS.n3960 VSS.n2215 48.7629
R6050 VSS.n2964 VSS.n2213 48.7629
R6051 VSS.n4527 VSS.n1890 48.7629
R6052 VSS.n3153 VSS.n2498 48.7629
R6053 VSS.n3385 VSS.n2463 48.7629
R6054 VSS.n2905 VSS.n2904 48.7629
R6055 VSS.n1964 VSS.n1962 48.7629
R6056 VSS.t15 VSS.t20 45.5776
R6057 VSS.n4259 VSS.t77 42.6154
R6058 VSS.n4272 VSS.t82 42.5927
R6059 VSS.n4260 VSS.t76 42.4377
R6060 VSS.n4273 VSS.t81 42.3691
R6061 VSS.n867 VSS.n863 40.8246
R6062 VSS.n4855 VSS.n4854 40.8246
R6063 VSS.n4851 VSS.n874 40.8246
R6064 VSS.n4849 VSS.n873 40.8246
R6065 VSS.n4848 VSS.n4847 40.8246
R6066 VSS.n878 VSS.n872 40.8246
R6067 VSS.n880 VSS.n876 40.8246
R6068 VSS.n882 VSS.n871 40.8246
R6069 VSS.n884 VSS.n877 40.8246
R6070 VSS.n4844 VSS.n870 40.8246
R6071 VSS.n4845 VSS.n869 40.8246
R6072 VSS.n161 VSS.n157 40.8246
R6073 VSS.n5376 VSS.n5375 40.8246
R6074 VSS.n5372 VSS.n168 40.8246
R6075 VSS.n5370 VSS.n167 40.8246
R6076 VSS.n5369 VSS.n5368 40.8246
R6077 VSS.n172 VSS.n166 40.8246
R6078 VSS.n174 VSS.n170 40.8246
R6079 VSS.n176 VSS.n165 40.8246
R6080 VSS.n178 VSS.n171 40.8246
R6081 VSS.n5365 VSS.n164 40.8246
R6082 VSS.n5366 VSS.n163 40.8246
R6083 VSS.n581 VSS.n574 40.8246
R6084 VSS.n606 VSS.n605 40.8246
R6085 VSS.n602 VSS.n582 40.8246
R6086 VSS.n600 VSS.n580 40.8246
R6087 VSS.n599 VSS.n598 40.8246
R6088 VSS.n586 VSS.n579 40.8246
R6089 VSS.n588 VSS.n584 40.8246
R6090 VSS.n590 VSS.n578 40.8246
R6091 VSS.n592 VSS.n585 40.8246
R6092 VSS.n595 VSS.n577 40.8246
R6093 VSS.n596 VSS.n575 40.8246
R6094 VSS.n5352 VSS.n196 40.8246
R6095 VSS.n5352 VSS.n5351 40.8246
R6096 VSS.n207 VSS.n204 40.8246
R6097 VSS.n207 VSS.n199 40.8246
R6098 VSS.n211 VSS.n205 40.8246
R6099 VSS.n211 VSS.n200 40.8246
R6100 VSS.n217 VSS.n216 40.8246
R6101 VSS.n216 VSS.n201 40.8246
R6102 VSS.n5348 VSS.n5347 40.8246
R6103 VSS.n5344 VSS.n198 40.8246
R6104 VSS.n196 VSS.n194 40.8246
R6105 VSS.n5347 VSS.n198 40.8246
R6106 VSS.n5349 VSS.n5348 40.8246
R6107 VSS.n202 VSS.n201 40.8246
R6108 VSS.n206 VSS.n200 40.8246
R6109 VSS.n217 VSS.n206 40.8246
R6110 VSS.n209 VSS.n199 40.8246
R6111 VSS.n209 VSS.n205 40.8246
R6112 VSS.n5351 VSS.n197 40.8246
R6113 VSS.n204 VSS.n197 40.8246
R6114 VSS.n3668 VSS.n3633 40.8246
R6115 VSS.n3667 VSS.n3666 40.8246
R6116 VSS.n3665 VSS.n3664 40.8246
R6117 VSS.n3661 VSS.n3637 40.8246
R6118 VSS.n3660 VSS.n3659 40.8246
R6119 VSS.n3658 VSS.n3657 40.8246
R6120 VSS.n3656 VSS.n3655 40.8246
R6121 VSS.n3652 VSS.n3640 40.8246
R6122 VSS.n3651 VSS.n3650 40.8246
R6123 VSS.n3649 VSS.n3648 40.8246
R6124 VSS.n3648 VSS.n3647 40.8246
R6125 VSS.n3645 VSS.n270 40.8246
R6126 VSS.n3650 VSS.n3649 40.8246
R6127 VSS.n3652 VSS.n3651 40.8246
R6128 VSS.n3655 VSS.n3640 40.8246
R6129 VSS.n3657 VSS.n3656 40.8246
R6130 VSS.n3659 VSS.n3658 40.8246
R6131 VSS.n3661 VSS.n3660 40.8246
R6132 VSS.n3664 VSS.n3637 40.8246
R6133 VSS.n3666 VSS.n3665 40.8246
R6134 VSS.n3668 VSS.n3667 40.8246
R6135 VSS.n3633 VSS.n220 40.8246
R6136 VSS.n4970 VSS.n4969 40.8246
R6137 VSS.n4982 VSS.n4971 40.8246
R6138 VSS.n4994 VSS.n4993 40.8246
R6139 VSS.n4990 VSS.n4972 40.8246
R6140 VSS.n4988 VSS.n4981 40.8246
R6141 VSS.n4986 VSS.n4973 40.8246
R6142 VSS.n4984 VSS.n4980 40.8246
R6143 VSS.n4979 VSS.n4974 40.8246
R6144 VSS.n4997 VSS.n4996 40.8246
R6145 VSS.n4999 VSS.n4975 40.8246
R6146 VSS.n4999 VSS.n4977 40.8246
R6147 VSS.n5003 VSS.n271 40.8246
R6148 VSS.n4997 VSS.n4975 40.8246
R6149 VSS.n4996 VSS.n4979 40.8246
R6150 VSS.n4984 VSS.n4974 40.8246
R6151 VSS.n4986 VSS.n4980 40.8246
R6152 VSS.n4988 VSS.n4973 40.8246
R6153 VSS.n4990 VSS.n4981 40.8246
R6154 VSS.n4993 VSS.n4972 40.8246
R6155 VSS.n4994 VSS.n4982 40.8246
R6156 VSS.n4971 VSS.n4970 40.8246
R6157 VSS.n5006 VSS.n4969 40.8246
R6158 VSS.n674 VSS.n671 40.8246
R6159 VSS.n5046 VSS.n5045 40.8246
R6160 VSS.n5042 VSS.n681 40.8246
R6161 VSS.n5040 VSS.n680 40.8246
R6162 VSS.n5039 VSS.n5038 40.8246
R6163 VSS.n685 VSS.n679 40.8246
R6164 VSS.n687 VSS.n683 40.8246
R6165 VSS.n689 VSS.n678 40.8246
R6166 VSS.n691 VSS.n684 40.8246
R6167 VSS.n5035 VSS.n677 40.8246
R6168 VSS.n5036 VSS.n676 40.8246
R6169 VSS.n705 VSS.n698 40.8246
R6170 VSS.n5025 VSS.n5024 40.8246
R6171 VSS.n5021 VSS.n706 40.8246
R6172 VSS.n5019 VSS.n704 40.8246
R6173 VSS.n5018 VSS.n5017 40.8246
R6174 VSS.n710 VSS.n703 40.8246
R6175 VSS.n712 VSS.n708 40.8246
R6176 VSS.n714 VSS.n702 40.8246
R6177 VSS.n716 VSS.n709 40.8246
R6178 VSS.n5014 VSS.n701 40.8246
R6179 VSS.n5015 VSS.n699 40.8246
R6180 VSS.n5015 VSS.n5014 40.8246
R6181 VSS.n716 VSS.n701 40.8246
R6182 VSS.n714 VSS.n709 40.8246
R6183 VSS.n712 VSS.n702 40.8246
R6184 VSS.n710 VSS.n708 40.8246
R6185 VSS.n5017 VSS.n703 40.8246
R6186 VSS.n5019 VSS.n5018 40.8246
R6187 VSS.n5021 VSS.n704 40.8246
R6188 VSS.n5024 VSS.n706 40.8246
R6189 VSS.n5025 VSS.n705 40.8246
R6190 VSS.n5027 VSS.n698 40.8246
R6191 VSS.n4196 VSS.n4195 40.8246
R6192 VSS.n4194 VSS.n4193 40.8246
R6193 VSS.n5449 VSS.n68 40.8246
R6194 VSS.n5448 VSS.n5447 40.8246
R6195 VSS.n5446 VSS.n5445 40.8246
R6196 VSS.n546 VSS.n72 40.8246
R6197 VSS.n548 VSS.n547 40.8246
R6198 VSS.n550 VSS.n549 40.8246
R6199 VSS.n562 VSS.n544 40.8246
R6200 VSS.n565 VSS.n563 40.8246
R6201 VSS.n565 VSS.n564 40.8246
R6202 VSS.n571 VSS.n570 40.8246
R6203 VSS.n569 VSS.n568 40.8246
R6204 VSS.n5154 VSS.n372 40.8246
R6205 VSS.n5153 VSS.n5152 40.8246
R6206 VSS.n3758 VSS.n373 40.8246
R6207 VSS.n3760 VSS.n3759 40.8246
R6208 VSS.n3767 VSS.n3756 40.8246
R6209 VSS.n3769 VSS.n3768 40.8246
R6210 VSS.n3776 VSS.n3752 40.8246
R6211 VSS.n3779 VSS.n3777 40.8246
R6212 VSS.n3778 VSS.n189 40.8246
R6213 VSS.n2266 VSS.n193 40.8246
R6214 VSS.n3878 VSS.n2259 40.8246
R6215 VSS.n3877 VSS.n3876 40.8246
R6216 VSS.n3875 VSS.n3874 40.8246
R6217 VSS.n3540 VSS.n2262 40.8246
R6218 VSS.n3546 VSS.n3541 40.8246
R6219 VSS.n3545 VSS.n3544 40.8246
R6220 VSS.n3543 VSS.n3542 40.8246
R6221 VSS.n3562 VSS.n2310 40.8246
R6222 VSS.n3565 VSS.n3563 40.8246
R6223 VSS.n3564 VSS.n693 40.8246
R6224 VSS.n754 VSS.n695 40.8246
R6225 VSS.n756 VSS.n755 40.8246
R6226 VSS.n4926 VSS.n757 40.8246
R6227 VSS.n4925 VSS.n4924 40.8246
R6228 VSS.n1130 VSS.n758 40.8246
R6229 VSS.n1132 VSS.n1131 40.8246
R6230 VSS.n1139 VSS.n1128 40.8246
R6231 VSS.n1141 VSS.n1140 40.8246
R6232 VSS.n1148 VSS.n1124 40.8246
R6233 VSS.n1151 VSS.n1149 40.8246
R6234 VSS.n1150 VSS.n886 40.8246
R6235 VSS.n4838 VSS.n4837 40.8246
R6236 VSS.n1299 VSS.n889 40.8246
R6237 VSS.n1610 VSS.n1300 40.8246
R6238 VSS.n1609 VSS.n1608 40.8246
R6239 VSS.n1607 VSS.n1606 40.8246
R6240 VSS.n1312 VSS.n1302 40.8246
R6241 VSS.n1595 VSS.n1313 40.8246
R6242 VSS.n1594 VSS.n1593 40.8246
R6243 VSS.n1592 VSS.n1591 40.8246
R6244 VSS.n1384 VSS.n1315 40.8246
R6245 VSS.n1385 VSS.n1384 40.8246
R6246 VSS.n4195 VSS.n4194 40.8246
R6247 VSS.n5449 VSS.n5448 40.8246
R6248 VSS.n5445 VSS.n72 40.8246
R6249 VSS.n549 VSS.n548 40.8246
R6250 VSS.n563 VSS.n562 40.8246
R6251 VSS.n568 VSS.n372 40.8246
R6252 VSS.n5152 VSS.n373 40.8246
R6253 VSS.n3760 VSS.n3756 40.8246
R6254 VSS.n3769 VSS.n3752 40.8246
R6255 VSS.n3779 VSS.n3778 40.8246
R6256 VSS.n5356 VSS.n193 40.8246
R6257 VSS.n3878 VSS.n3877 40.8246
R6258 VSS.n3874 VSS.n2262 40.8246
R6259 VSS.n3546 VSS.n3545 40.8246
R6260 VSS.n3542 VSS.n2310 40.8246
R6261 VSS.n3565 VSS.n3564 40.8246
R6262 VSS.n5030 VSS.n695 40.8246
R6263 VSS.n757 VSS.n756 40.8246
R6264 VSS.n4924 VSS.n758 40.8246
R6265 VSS.n1132 VSS.n1128 40.8246
R6266 VSS.n1141 VSS.n1124 40.8246
R6267 VSS.n1151 VSS.n1150 40.8246
R6268 VSS.n4837 VSS.n889 40.8246
R6269 VSS.n1610 VSS.n1609 40.8246
R6270 VSS.n1606 VSS.n1302 40.8246
R6271 VSS.n1595 VSS.n1594 40.8246
R6272 VSS.n1591 VSS.n1315 40.8246
R6273 VSS.n1593 VSS.n1592 40.8246
R6274 VSS.n1313 VSS.n1312 40.8246
R6275 VSS.n1608 VSS.n1607 40.8246
R6276 VSS.n1300 VSS.n1299 40.8246
R6277 VSS.n4839 VSS.n4838 40.8246
R6278 VSS.n1149 VSS.n1148 40.8246
R6279 VSS.n1140 VSS.n1139 40.8246
R6280 VSS.n1131 VSS.n1130 40.8246
R6281 VSS.n4926 VSS.n4925 40.8246
R6282 VSS.n755 VSS.n754 40.8246
R6283 VSS.n3563 VSS.n3562 40.8246
R6284 VSS.n3544 VSS.n3543 40.8246
R6285 VSS.n3541 VSS.n3540 40.8246
R6286 VSS.n3876 VSS.n3875 40.8246
R6287 VSS.n2266 VSS.n2259 40.8246
R6288 VSS.n3777 VSS.n3776 40.8246
R6289 VSS.n3768 VSS.n3767 40.8246
R6290 VSS.n3759 VSS.n3758 40.8246
R6291 VSS.n5154 VSS.n5153 40.8246
R6292 VSS.n570 VSS.n569 40.8246
R6293 VSS.n550 VSS.n544 40.8246
R6294 VSS.n547 VSS.n546 40.8246
R6295 VSS.n5447 VSS.n5446 40.8246
R6296 VSS.n4193 VSS.n68 40.8246
R6297 VSS.n4197 VSS.n4196 40.8246
R6298 VSS.n991 VSS.n967 40.8246
R6299 VSS.n989 VSS.n965 40.8246
R6300 VSS.n988 VSS.n987 40.8246
R6301 VSS.n972 VSS.n964 40.8246
R6302 VSS.n974 VSS.n969 40.8246
R6303 VSS.n976 VSS.n963 40.8246
R6304 VSS.n978 VSS.n970 40.8246
R6305 VSS.n971 VSS.n962 40.8246
R6306 VSS.n985 VSS.n984 40.8246
R6307 VSS.n981 VSS.n961 40.8246
R6308 VSS.n996 VSS.n957 40.8246
R6309 VSS.n981 VSS.n957 40.8246
R6310 VSS.n984 VSS.n961 40.8246
R6311 VSS.n985 VSS.n971 40.8246
R6312 VSS.n978 VSS.n962 40.8246
R6313 VSS.n976 VSS.n970 40.8246
R6314 VSS.n974 VSS.n963 40.8246
R6315 VSS.n972 VSS.n969 40.8246
R6316 VSS.n987 VSS.n964 40.8246
R6317 VSS.n989 VSS.n988 40.8246
R6318 VSS.n991 VSS.n965 40.8246
R6319 VSS.n994 VSS.n967 40.8246
R6320 VSS.n1032 VSS.n1031 40.8246
R6321 VSS.n1030 VSS.n1029 40.8246
R6322 VSS.n1028 VSS.n1027 40.8246
R6323 VSS.n1024 VSS.n1001 40.8246
R6324 VSS.n1023 VSS.n1022 40.8246
R6325 VSS.n1021 VSS.n1020 40.8246
R6326 VSS.n1019 VSS.n1018 40.8246
R6327 VSS.n1015 VSS.n1004 40.8246
R6328 VSS.n1014 VSS.n1013 40.8246
R6329 VSS.n1012 VSS.n1011 40.8246
R6330 VSS.n1011 VSS.n1007 40.8246
R6331 VSS.n5328 VSS.n272 40.8246
R6332 VSS.n1013 VSS.n1012 40.8246
R6333 VSS.n1015 VSS.n1014 40.8246
R6334 VSS.n1018 VSS.n1004 40.8246
R6335 VSS.n1020 VSS.n1019 40.8246
R6336 VSS.n1022 VSS.n1021 40.8246
R6337 VSS.n1024 VSS.n1023 40.8246
R6338 VSS.n1027 VSS.n1001 40.8246
R6339 VSS.n1029 VSS.n1028 40.8246
R6340 VSS.n1031 VSS.n1030 40.8246
R6341 VSS.n1033 VSS.n1032 40.8246
R6342 VSS.n4096 VSS.n4095 40.8246
R6343 VSS.n4094 VSS.n4093 40.8246
R6344 VSS.n5470 VSS.n26 40.8246
R6345 VSS.n5469 VSS.n5468 40.8246
R6346 VSS.n5467 VSS.n5466 40.8246
R6347 VSS.n465 VSS.n30 40.8246
R6348 VSS.n467 VSS.n466 40.8246
R6349 VSS.n469 VSS.n468 40.8246
R6350 VSS.n519 VSS.n460 40.8246
R6351 VSS.n522 VSS.n520 40.8246
R6352 VSS.n522 VSS.n521 40.8246
R6353 VSS.n5174 VSS.n232 40.8246
R6354 VSS.n5173 VSS.n5172 40.8246
R6355 VSS.n3677 VSS.n338 40.8246
R6356 VSS.n3679 VSS.n3678 40.8246
R6357 VSS.n3681 VSS.n3680 40.8246
R6358 VSS.n3695 VSS.n3676 40.8246
R6359 VSS.n3697 VSS.n3696 40.8246
R6360 VSS.n3701 VSS.n3698 40.8246
R6361 VSS.n3700 VSS.n3699 40.8246
R6362 VSS.n3803 VSS.n3671 40.8246
R6363 VSS.n3805 VSS.n3804 40.8246
R6364 VSS.n3809 VSS.n3808 40.8246
R6365 VSS.n3843 VSS.n2277 40.8246
R6366 VSS.n3842 VSS.n3841 40.8246
R6367 VSS.n3840 VSS.n3839 40.8246
R6368 VSS.n2288 VSS.n2280 40.8246
R6369 VSS.n2291 VSS.n2289 40.8246
R6370 VSS.n3618 VSS.n2292 40.8246
R6371 VSS.n3617 VSS.n3616 40.8246
R6372 VSS.n2298 VSS.n2293 40.8246
R6373 VSS.n2301 VSS.n2299 40.8246
R6374 VSS.n2300 VSS.n718 40.8246
R6375 VSS.n4966 VSS.n4965 40.8246
R6376 VSS.n4964 VSS.n4963 40.8246
R6377 VSS.n1047 VSS.n721 40.8246
R6378 VSS.n1056 VSS.n1046 40.8246
R6379 VSS.n1058 VSS.n1057 40.8246
R6380 VSS.n1062 VSS.n1059 40.8246
R6381 VSS.n1061 VSS.n1060 40.8246
R6382 VSS.n1080 VSS.n1040 40.8246
R6383 VSS.n1082 VSS.n1081 40.8246
R6384 VSS.n1175 VSS.n1035 40.8246
R6385 VSS.n1177 VSS.n1176 40.8246
R6386 VSS.n1181 VSS.n1180 40.8246
R6387 VSS.n4828 VSS.n914 40.8246
R6388 VSS.n4827 VSS.n4826 40.8246
R6389 VSS.n1354 VSS.n915 40.8246
R6390 VSS.n1361 VSS.n1353 40.8246
R6391 VSS.n1363 VSS.n1362 40.8246
R6392 VSS.n1370 VSS.n1347 40.8246
R6393 VSS.n1372 VSS.n1371 40.8246
R6394 VSS.n1379 VSS.n1343 40.8246
R6395 VSS.n1559 VSS.n1380 40.8246
R6396 VSS.n1559 VSS.n1558 40.8246
R6397 VSS.n4095 VSS.n4094 40.8246
R6398 VSS.n5470 VSS.n5469 40.8246
R6399 VSS.n5466 VSS.n30 40.8246
R6400 VSS.n468 VSS.n467 40.8246
R6401 VSS.n520 VSS.n519 40.8246
R6402 VSS.n5172 VSS.n338 40.8246
R6403 VSS.n3680 VSS.n3679 40.8246
R6404 VSS.n3696 VSS.n3695 40.8246
R6405 VSS.n3701 VSS.n3700 40.8246
R6406 VSS.n3804 VSS.n3803 40.8246
R6407 VSS.n3808 VSS.n222 40.8246
R6408 VSS.n3843 VSS.n3842 40.8246
R6409 VSS.n3839 VSS.n2280 40.8246
R6410 VSS.n2292 VSS.n2291 40.8246
R6411 VSS.n3616 VSS.n2293 40.8246
R6412 VSS.n2301 VSS.n2300 40.8246
R6413 VSS.n5009 VSS.n4966 40.8246
R6414 VSS.n4963 VSS.n721 40.8246
R6415 VSS.n1057 VSS.n1056 40.8246
R6416 VSS.n1062 VSS.n1061 40.8246
R6417 VSS.n1081 VSS.n1080 40.8246
R6418 VSS.n1176 VSS.n1175 40.8246
R6419 VSS.n1181 VSS.n914 40.8246
R6420 VSS.n4826 VSS.n915 40.8246
R6421 VSS.n1362 VSS.n1361 40.8246
R6422 VSS.n1371 VSS.n1370 40.8246
R6423 VSS.n1380 VSS.n1379 40.8246
R6424 VSS.n1372 VSS.n1343 40.8246
R6425 VSS.n1363 VSS.n1347 40.8246
R6426 VSS.n1354 VSS.n1353 40.8246
R6427 VSS.n4828 VSS.n4827 40.8246
R6428 VSS.n1180 VSS.n1179 40.8246
R6429 VSS.n1082 VSS.n1035 40.8246
R6430 VSS.n1060 VSS.n1040 40.8246
R6431 VSS.n1059 VSS.n1058 40.8246
R6432 VSS.n1047 VSS.n1046 40.8246
R6433 VSS.n4965 VSS.n4964 40.8246
R6434 VSS.n2299 VSS.n2298 40.8246
R6435 VSS.n3618 VSS.n3617 40.8246
R6436 VSS.n2289 VSS.n2288 40.8246
R6437 VSS.n3841 VSS.n3840 40.8246
R6438 VSS.n3809 VSS.n2277 40.8246
R6439 VSS.n3699 VSS.n3671 40.8246
R6440 VSS.n3698 VSS.n3697 40.8246
R6441 VSS.n3681 VSS.n3676 40.8246
R6442 VSS.n3678 VSS.n3677 40.8246
R6443 VSS.n5174 VSS.n5173 40.8246
R6444 VSS.n469 VSS.n460 40.8246
R6445 VSS.n466 VSS.n465 40.8246
R6446 VSS.n5468 VSS.n5467 40.8246
R6447 VSS.n4093 VSS.n26 40.8246
R6448 VSS.n4097 VSS.n4096 40.8246
R6449 VSS.n235 VSS.n234 40.8246
R6450 VSS.n248 VSS.n236 40.8246
R6451 VSS.n260 VSS.n259 40.8246
R6452 VSS.n256 VSS.n237 40.8246
R6453 VSS.n254 VSS.n247 40.8246
R6454 VSS.n252 VSS.n238 40.8246
R6455 VSS.n250 VSS.n246 40.8246
R6456 VSS.n245 VSS.n239 40.8246
R6457 VSS.n263 VSS.n262 40.8246
R6458 VSS.n265 VSS.n240 40.8246
R6459 VSS.n265 VSS.n242 40.8246
R6460 VSS.n5330 VSS.n243 40.8246
R6461 VSS.n263 VSS.n240 40.8246
R6462 VSS.n262 VSS.n245 40.8246
R6463 VSS.n250 VSS.n239 40.8246
R6464 VSS.n252 VSS.n246 40.8246
R6465 VSS.n254 VSS.n238 40.8246
R6466 VSS.n256 VSS.n247 40.8246
R6467 VSS.n259 VSS.n237 40.8246
R6468 VSS.n260 VSS.n248 40.8246
R6469 VSS.n5337 VSS.n232 40.8246
R6470 VSS.n521 VSS.n228 40.8246
R6471 VSS.n236 VSS.n235 40.8246
R6472 VSS.n5334 VSS.n234 40.8246
R6473 VSS.n596 VSS.n595 40.8246
R6474 VSS.n592 VSS.n577 40.8246
R6475 VSS.n590 VSS.n585 40.8246
R6476 VSS.n588 VSS.n578 40.8246
R6477 VSS.n586 VSS.n584 40.8246
R6478 VSS.n598 VSS.n579 40.8246
R6479 VSS.n600 VSS.n599 40.8246
R6480 VSS.n602 VSS.n580 40.8246
R6481 VSS.n605 VSS.n582 40.8246
R6482 VSS.n606 VSS.n581 40.8246
R6483 VSS.n572 VSS.n571 40.8246
R6484 VSS.n564 VSS.n182 40.8246
R6485 VSS.n608 VSS.n574 40.8246
R6486 VSS.n5366 VSS.n5365 40.8246
R6487 VSS.n178 VSS.n164 40.8246
R6488 VSS.n176 VSS.n171 40.8246
R6489 VSS.n174 VSS.n165 40.8246
R6490 VSS.n172 VSS.n170 40.8246
R6491 VSS.n5368 VSS.n166 40.8246
R6492 VSS.n5370 VSS.n5369 40.8246
R6493 VSS.n5372 VSS.n167 40.8246
R6494 VSS.n5375 VSS.n168 40.8246
R6495 VSS.n5036 VSS.n5035 40.8246
R6496 VSS.n691 VSS.n677 40.8246
R6497 VSS.n689 VSS.n684 40.8246
R6498 VSS.n687 VSS.n678 40.8246
R6499 VSS.n685 VSS.n683 40.8246
R6500 VSS.n5038 VSS.n679 40.8246
R6501 VSS.n5040 VSS.n5039 40.8246
R6502 VSS.n5042 VSS.n680 40.8246
R6503 VSS.n5045 VSS.n681 40.8246
R6504 VSS.n4845 VSS.n4844 40.8246
R6505 VSS.n884 VSS.n870 40.8246
R6506 VSS.n882 VSS.n877 40.8246
R6507 VSS.n880 VSS.n871 40.8246
R6508 VSS.n878 VSS.n876 40.8246
R6509 VSS.n4847 VSS.n872 40.8246
R6510 VSS.n4849 VSS.n4848 40.8246
R6511 VSS.n4851 VSS.n873 40.8246
R6512 VSS.n4854 VSS.n874 40.8246
R6513 VSS.n2185 VSS.n2173 40.8246
R6514 VSS.n2184 VSS.n2174 40.8246
R6515 VSS.n2196 VSS.n2195 40.8246
R6516 VSS.n2192 VSS.n2175 40.8246
R6517 VSS.n2190 VSS.n2183 40.8246
R6518 VSS.n2188 VSS.n2176 40.8246
R6519 VSS.n2182 VSS.n2181 40.8246
R6520 VSS.n2199 VSS.n2177 40.8246
R6521 VSS.n2198 VSS.n2178 40.8246
R6522 VSS.n2204 VSS.n2203 40.8246
R6523 VSS.n2203 VSS.n2179 40.8246
R6524 VSS.n3155 VSS.n2495 40.8246
R6525 VSS.n2204 VSS.n2178 40.8246
R6526 VSS.n2199 VSS.n2198 40.8246
R6527 VSS.n2181 VSS.n2177 40.8246
R6528 VSS.n2188 VSS.n2182 40.8246
R6529 VSS.n2190 VSS.n2176 40.8246
R6530 VSS.n2192 VSS.n2183 40.8246
R6531 VSS.n2195 VSS.n2175 40.8246
R6532 VSS.n2196 VSS.n2184 40.8246
R6533 VSS.n2185 VSS.n2174 40.8246
R6534 VSS.n2206 VSS.n2173 40.8246
R6535 VSS.n3419 VSS.n3387 40.8246
R6536 VSS.n3398 VSS.n3388 40.8246
R6537 VSS.n3398 VSS.n3394 40.8246
R6538 VSS.n3402 VSS.n3389 40.8246
R6539 VSS.n3402 VSS.n3395 40.8246
R6540 VSS.n3406 VSS.n3390 40.8246
R6541 VSS.n3406 VSS.n3396 40.8246
R6542 VSS.n3397 VSS.n3391 40.8246
R6543 VSS.n3414 VSS.n3397 40.8246
R6544 VSS.n3393 VSS.n3392 40.8246
R6545 VSS.n3417 VSS.n3416 40.8246
R6546 VSS.n3416 VSS.n3393 40.8246
R6547 VSS.n3414 VSS.n3413 40.8246
R6548 VSS.n3413 VSS.n3392 40.8246
R6549 VSS.n3408 VSS.n3396 40.8246
R6550 VSS.n3408 VSS.n3391 40.8246
R6551 VSS.n3404 VSS.n3395 40.8246
R6552 VSS.n3404 VSS.n3390 40.8246
R6553 VSS.n3400 VSS.n3394 40.8246
R6554 VSS.n3400 VSS.n3389 40.8246
R6555 VSS.n3953 VSS.n3952 40.8246
R6556 VSS.n3951 VSS.n3950 40.8246
R6557 VSS.n3949 VSS.n3948 40.8246
R6558 VSS.n3945 VSS.n3925 40.8246
R6559 VSS.n3944 VSS.n3943 40.8246
R6560 VSS.n3942 VSS.n3941 40.8246
R6561 VSS.n3940 VSS.n3939 40.8246
R6562 VSS.n3936 VSS.n3928 40.8246
R6563 VSS.n3935 VSS.n3934 40.8246
R6564 VSS.n3933 VSS.n3932 40.8246
R6565 VSS.n3932 VSS.n3931 40.8246
R6566 VSS.n3934 VSS.n3933 40.8246
R6567 VSS.n3936 VSS.n3935 40.8246
R6568 VSS.n3939 VSS.n3928 40.8246
R6569 VSS.n3941 VSS.n3940 40.8246
R6570 VSS.n3943 VSS.n3942 40.8246
R6571 VSS.n3945 VSS.n3944 40.8246
R6572 VSS.n3948 VSS.n3925 40.8246
R6573 VSS.n3950 VSS.n3949 40.8246
R6574 VSS.n3952 VSS.n3951 40.8246
R6575 VSS.n3954 VSS.n3953 40.8246
R6576 VSS.n661 VSS.n657 40.8246
R6577 VSS.n5083 VSS.n5082 40.8246
R6578 VSS.n5079 VSS.n5059 40.8246
R6579 VSS.n5077 VSS.n5058 40.8246
R6580 VSS.n5076 VSS.n5075 40.8246
R6581 VSS.n5063 VSS.n5057 40.8246
R6582 VSS.n5065 VSS.n5061 40.8246
R6583 VSS.n5067 VSS.n5056 40.8246
R6584 VSS.n5069 VSS.n5062 40.8246
R6585 VSS.n5072 VSS.n5055 40.8246
R6586 VSS.n5073 VSS.n5054 40.8246
R6587 VSS.n5073 VSS.n5072 40.8246
R6588 VSS.n5069 VSS.n5055 40.8246
R6589 VSS.n5067 VSS.n5062 40.8246
R6590 VSS.n5065 VSS.n5056 40.8246
R6591 VSS.n5063 VSS.n5061 40.8246
R6592 VSS.n5075 VSS.n5057 40.8246
R6593 VSS.n5077 VSS.n5076 40.8246
R6594 VSS.n5079 VSS.n5058 40.8246
R6595 VSS.n5082 VSS.n5059 40.8246
R6596 VSS.n5412 VSS.n5411 40.8246
R6597 VSS.n5410 VSS.n5409 40.8246
R6598 VSS.n5408 VSS.n5407 40.8246
R6599 VSS.n136 VSS.n131 40.8246
R6600 VSS.n138 VSS.n137 40.8246
R6601 VSS.n5396 VSS.n139 40.8246
R6602 VSS.n5395 VSS.n5394 40.8246
R6603 VSS.n152 VSS.n140 40.8246
R6604 VSS.n154 VSS.n153 40.8246
R6605 VSS.n5383 VSS.n155 40.8246
R6606 VSS.n5382 VSS.n5381 40.8246
R6607 VSS.n5119 VSS.n5118 40.8246
R6608 VSS.n5117 VSS.n5116 40.8246
R6609 VSS.n5115 VSS.n5114 40.8246
R6610 VSS.n636 VSS.n631 40.8246
R6611 VSS.n638 VSS.n637 40.8246
R6612 VSS.n5103 VSS.n639 40.8246
R6613 VSS.n5102 VSS.n5101 40.8246
R6614 VSS.n652 VSS.n640 40.8246
R6615 VSS.n654 VSS.n653 40.8246
R6616 VSS.n5090 VSS.n655 40.8246
R6617 VSS.n5089 VSS.n5088 40.8246
R6618 VSS.n2421 VSS.n2420 40.8246
R6619 VSS.n3908 VSS.n2245 40.8246
R6620 VSS.n3907 VSS.n3906 40.8246
R6621 VSS.n3475 VSS.n2246 40.8246
R6622 VSS.n3477 VSS.n3476 40.8246
R6623 VSS.n3484 VSS.n3471 40.8246
R6624 VSS.n3488 VSS.n3485 40.8246
R6625 VSS.n3487 VSS.n3486 40.8246
R6626 VSS.n3506 VSS.n3466 40.8246
R6627 VSS.n3509 VSS.n3507 40.8246
R6628 VSS.n3508 VSS.n668 40.8246
R6629 VSS.n4891 VSS.n4890 40.8246
R6630 VSS.n4889 VSS.n4888 40.8246
R6631 VSS.n4887 VSS.n4886 40.8246
R6632 VSS.n843 VSS.n838 40.8246
R6633 VSS.n845 VSS.n844 40.8246
R6634 VSS.n4875 VSS.n846 40.8246
R6635 VSS.n4874 VSS.n4873 40.8246
R6636 VSS.n859 VSS.n847 40.8246
R6637 VSS.n861 VSS.n860 40.8246
R6638 VSS.n4862 VSS.n862 40.8246
R6639 VSS.n4861 VSS.n4860 40.8246
R6640 VSS.n4741 VSS.n4740 40.8246
R6641 VSS.n4770 VSS.n1278 40.8246
R6642 VSS.n4769 VSS.n4768 40.8246
R6643 VSS.n1416 VSS.n1279 40.8246
R6644 VSS.n1423 VSS.n1415 40.8246
R6645 VSS.n1431 VSS.n1424 40.8246
R6646 VSS.n1430 VSS.n1429 40.8246
R6647 VSS.n1428 VSS.n1427 40.8246
R6648 VSS.n1426 VSS.n1425 40.8246
R6649 VSS.n1482 VSS.n1409 40.8246
R6650 VSS.n1484 VSS.n1483 40.8246
R6651 VSS.n4529 VSS.n4528 40.8246
R6652 VSS.n4540 VSS.n4530 40.8246
R6653 VSS.n4550 VSS.n4549 40.8246
R6654 VSS.n4546 VSS.n4531 40.8246
R6655 VSS.n4544 VSS.n4539 40.8246
R6656 VSS.n4542 VSS.n4532 40.8246
R6657 VSS.n4538 VSS.n4537 40.8246
R6658 VSS.n4553 VSS.n4533 40.8246
R6659 VSS.n4552 VSS.n4534 40.8246
R6660 VSS.n4558 VSS.n4557 40.8246
R6661 VSS.n4557 VSS.n4535 40.8246
R6662 VSS.n4558 VSS.n4534 40.8246
R6663 VSS.n4553 VSS.n4552 40.8246
R6664 VSS.n4537 VSS.n4533 40.8246
R6665 VSS.n4542 VSS.n4538 40.8246
R6666 VSS.n4544 VSS.n4532 40.8246
R6667 VSS.n4546 VSS.n4539 40.8246
R6668 VSS.n4549 VSS.n4531 40.8246
R6669 VSS.n4550 VSS.n4540 40.8246
R6670 VSS.n4530 VSS.n4529 40.8246
R6671 VSS.n4560 VSS.n4528 40.8246
R6672 VSS.n2929 VSS.n2907 40.8246
R6673 VSS.n2997 VSS.n2996 40.8246
R6674 VSS.n2993 VSS.n2971 40.8246
R6675 VSS.n2991 VSS.n2970 40.8246
R6676 VSS.n2990 VSS.n2989 40.8246
R6677 VSS.n2975 VSS.n2969 40.8246
R6678 VSS.n2977 VSS.n2973 40.8246
R6679 VSS.n2979 VSS.n2968 40.8246
R6680 VSS.n2981 VSS.n2974 40.8246
R6681 VSS.n2986 VSS.n2967 40.8246
R6682 VSS.n2987 VSS.n2965 40.8246
R6683 VSS.n2987 VSS.n2986 40.8246
R6684 VSS.n2981 VSS.n2967 40.8246
R6685 VSS.n2979 VSS.n2974 40.8246
R6686 VSS.n2977 VSS.n2968 40.8246
R6687 VSS.n2975 VSS.n2973 40.8246
R6688 VSS.n2989 VSS.n2969 40.8246
R6689 VSS.n2991 VSS.n2990 40.8246
R6690 VSS.n2993 VSS.n2970 40.8246
R6691 VSS.n2996 VSS.n2971 40.8246
R6692 VSS.n2962 VSS.n2961 40.8246
R6693 VSS.n2958 VSS.n2932 40.8246
R6694 VSS.n2957 VSS.n2956 40.8246
R6695 VSS.n2955 VSS.n2954 40.8246
R6696 VSS.n2953 VSS.n2952 40.8246
R6697 VSS.n2949 VSS.n2935 40.8246
R6698 VSS.n2948 VSS.n2947 40.8246
R6699 VSS.n2946 VSS.n2945 40.8246
R6700 VSS.n2944 VSS.n2943 40.8246
R6701 VSS.n2940 VSS.n2938 40.8246
R6702 VSS.n2940 VSS.n2939 40.8246
R6703 VSS.n2943 VSS.n2938 40.8246
R6704 VSS.n2945 VSS.n2944 40.8246
R6705 VSS.n2947 VSS.n2946 40.8246
R6706 VSS.n2949 VSS.n2948 40.8246
R6707 VSS.n2952 VSS.n2935 40.8246
R6708 VSS.n2954 VSS.n2953 40.8246
R6709 VSS.n2956 VSS.n2955 40.8246
R6710 VSS.n2958 VSS.n2957 40.8246
R6711 VSS.n2961 VSS.n2932 40.8246
R6712 VSS.n2963 VSS.n2962 40.8246
R6713 VSS.n3996 VSS.n2118 40.8246
R6714 VSS.n3995 VSS.n3994 40.8246
R6715 VSS.n2130 VSS.n2119 40.8246
R6716 VSS.n2132 VSS.n2131 40.8246
R6717 VSS.n3983 VSS.n2133 40.8246
R6718 VSS.n3982 VSS.n3981 40.8246
R6719 VSS.n2142 VSS.n2134 40.8246
R6720 VSS.n3972 VSS.n2143 40.8246
R6721 VSS.n3971 VSS.n3970 40.8246
R6722 VSS.n3969 VSS.n3968 40.8246
R6723 VSS.n3963 VSS.n2146 40.8246
R6724 VSS.n3205 VSS.n3203 40.8246
R6725 VSS.n3342 VSS.n3206 40.8246
R6726 VSS.n3341 VSS.n3340 40.8246
R6727 VSS.n3339 VSS.n3338 40.8246
R6728 VSS.n3221 VSS.n3209 40.8246
R6729 VSS.n3224 VSS.n3222 40.8246
R6730 VSS.n3323 VSS.n3225 40.8246
R6731 VSS.n3322 VSS.n3321 40.8246
R6732 VSS.n3309 VSS.n3226 40.8246
R6733 VSS.n3312 VSS.n3310 40.8246
R6734 VSS.n3311 VSS.n2214 40.8246
R6735 VSS.n3920 VSS.n3919 40.8246
R6736 VSS.n3918 VSS.n3917 40.8246
R6737 VSS.n2354 VSS.n2219 40.8246
R6738 VSS.n2356 VSS.n2355 40.8246
R6739 VSS.n2363 VSS.n2345 40.8246
R6740 VSS.n2365 VSS.n2364 40.8246
R6741 VSS.n2372 VSS.n2344 40.8246
R6742 VSS.n2374 VSS.n2373 40.8246
R6743 VSS.n3439 VSS.n2331 40.8246
R6744 VSS.n3441 VSS.n3440 40.8246
R6745 VSS.n3443 VSS.n3442 40.8246
R6746 VSS.n2328 VSS.n2327 40.8246
R6747 VSS.n4595 VSS.n1840 40.8246
R6748 VSS.n4594 VSS.n4593 40.8246
R6749 VSS.n4592 VSS.n4591 40.8246
R6750 VSS.n1857 VSS.n1845 40.8246
R6751 VSS.n1860 VSS.n1858 40.8246
R6752 VSS.n4576 VSS.n1861 40.8246
R6753 VSS.n4575 VSS.n4574 40.8246
R6754 VSS.n1887 VSS.n1862 40.8246
R6755 VSS.n4565 VSS.n1888 40.8246
R6756 VSS.n4564 VSS.n4563 40.8246
R6757 VSS.n1949 VSS.n1948 40.8246
R6758 VSS.n1947 VSS.n1946 40.8246
R6759 VSS.n1945 VSS.n1944 40.8246
R6760 VSS.n1943 VSS.n1942 40.8246
R6761 VSS.n1903 VSS.n1893 40.8246
R6762 VSS.n1932 VSS.n1904 40.8246
R6763 VSS.n1931 VSS.n1930 40.8246
R6764 VSS.n1929 VSS.n1928 40.8246
R6765 VSS.n1918 VSS.n1906 40.8246
R6766 VSS.n1917 VSS.n1916 40.8246
R6767 VSS.n1915 VSS.n1250 40.8246
R6768 VSS.n2118 VSS.n2067 40.8246
R6769 VSS.n3994 VSS.n2119 40.8246
R6770 VSS.n2133 VSS.n2132 40.8246
R6771 VSS.n3981 VSS.n2134 40.8246
R6772 VSS.n3972 VSS.n3971 40.8246
R6773 VSS.n3968 VSS.n2146 40.8246
R6774 VSS.n3203 VSS.n2171 40.8246
R6775 VSS.n3342 VSS.n3341 40.8246
R6776 VSS.n3338 VSS.n3209 40.8246
R6777 VSS.n3225 VSS.n3224 40.8246
R6778 VSS.n3321 VSS.n3226 40.8246
R6779 VSS.n3312 VSS.n3311 40.8246
R6780 VSS.n3957 VSS.n3920 40.8246
R6781 VSS.n3917 VSS.n2219 40.8246
R6782 VSS.n2356 VSS.n2345 40.8246
R6783 VSS.n2365 VSS.n2344 40.8246
R6784 VSS.n2374 VSS.n2331 40.8246
R6785 VSS.n3442 VSS.n3441 40.8246
R6786 VSS.n2329 VSS.n2328 40.8246
R6787 VSS.n4595 VSS.n4594 40.8246
R6788 VSS.n4591 VSS.n1845 40.8246
R6789 VSS.n1861 VSS.n1860 40.8246
R6790 VSS.n4574 VSS.n1862 40.8246
R6791 VSS.n4565 VSS.n4564 40.8246
R6792 VSS.n1950 VSS.n1949 40.8246
R6793 VSS.n1888 VSS.n1887 40.8246
R6794 VSS.n4576 VSS.n4575 40.8246
R6795 VSS.n1858 VSS.n1857 40.8246
R6796 VSS.n4593 VSS.n4592 40.8246
R6797 VSS.n2327 VSS.n1840 40.8246
R6798 VSS.n3440 VSS.n3439 40.8246
R6799 VSS.n2373 VSS.n2372 40.8246
R6800 VSS.n2364 VSS.n2363 40.8246
R6801 VSS.n2355 VSS.n2354 40.8246
R6802 VSS.n3919 VSS.n3918 40.8246
R6803 VSS.n3310 VSS.n3309 40.8246
R6804 VSS.n3323 VSS.n3322 40.8246
R6805 VSS.n3222 VSS.n3221 40.8246
R6806 VSS.n3340 VSS.n3339 40.8246
R6807 VSS.n3206 VSS.n3205 40.8246
R6808 VSS.n3970 VSS.n3969 40.8246
R6809 VSS.n2143 VSS.n2142 40.8246
R6810 VSS.n3983 VSS.n3982 40.8246
R6811 VSS.n2131 VSS.n2130 40.8246
R6812 VSS.n3996 VSS.n3995 40.8246
R6813 VSS.n3060 VSS.n2778 40.8246
R6814 VSS.n2775 VSS.n2750 40.8246
R6815 VSS.n2775 VSS.n2774 40.8246
R6816 VSS.n2772 VSS.n2771 40.8246
R6817 VSS.n2771 VSS.n2751 40.8246
R6818 VSS.n2767 VSS.n2766 40.8246
R6819 VSS.n2766 VSS.n2765 40.8246
R6820 VSS.n2763 VSS.n2762 40.8246
R6821 VSS.n2762 VSS.n2754 40.8246
R6822 VSS.n2758 VSS.n2757 40.8246
R6823 VSS.n2756 VSS.n2461 40.8246
R6824 VSS.n2757 VSS.n2756 40.8246
R6825 VSS.n2759 VSS.n2754 40.8246
R6826 VSS.n2759 VSS.n2758 40.8246
R6827 VSS.n2765 VSS.n2764 40.8246
R6828 VSS.n2764 VSS.n2763 40.8246
R6829 VSS.n2768 VSS.n2751 40.8246
R6830 VSS.n2768 VSS.n2767 40.8246
R6831 VSS.n2774 VSS.n2773 40.8246
R6832 VSS.n2773 VSS.n2772 40.8246
R6833 VSS.n3025 VSS.n3024 40.8246
R6834 VSS.n3021 VSS.n2812 40.8246
R6835 VSS.n3021 VSS.n3020 40.8246
R6836 VSS.n3018 VSS.n3017 40.8246
R6837 VSS.n3017 VSS.n2813 40.8246
R6838 VSS.n3013 VSS.n3012 40.8246
R6839 VSS.n3012 VSS.n3011 40.8246
R6840 VSS.n3009 VSS.n3008 40.8246
R6841 VSS.n3008 VSS.n2816 40.8246
R6842 VSS.n3004 VSS.n3003 40.8246
R6843 VSS.n3002 VSS.n3001 40.8246
R6844 VSS.n3003 VSS.n3002 40.8246
R6845 VSS.n3005 VSS.n2816 40.8246
R6846 VSS.n3005 VSS.n3004 40.8246
R6847 VSS.n3011 VSS.n3010 40.8246
R6848 VSS.n3010 VSS.n3009 40.8246
R6849 VSS.n3014 VSS.n2813 40.8246
R6850 VSS.n3014 VSS.n3013 40.8246
R6851 VSS.n3020 VSS.n3019 40.8246
R6852 VSS.n3019 VSS.n3018 40.8246
R6853 VSS.n4496 VSS.n1997 40.8246
R6854 VSS.n4500 VSS.n4499 40.8246
R6855 VSS.n4501 VSS.n4500 40.8246
R6856 VSS.n4505 VSS.n1995 40.8246
R6857 VSS.n4506 VSS.n4505 40.8246
R6858 VSS.n4509 VSS.n4508 40.8246
R6859 VSS.n4509 VSS.n1993 40.8246
R6860 VSS.n4514 VSS.n4513 40.8246
R6861 VSS.n4515 VSS.n4514 40.8246
R6862 VSS.n4519 VSS.n1991 40.8246
R6863 VSS.n4521 VSS.n4520 40.8246
R6864 VSS.n4520 VSS.n4519 40.8246
R6865 VSS.n4516 VSS.n4515 40.8246
R6866 VSS.n4516 VSS.n1991 40.8246
R6867 VSS.n4512 VSS.n1993 40.8246
R6868 VSS.n4513 VSS.n4512 40.8246
R6869 VSS.n4507 VSS.n4506 40.8246
R6870 VSS.n4508 VSS.n4507 40.8246
R6871 VSS.n4502 VSS.n4501 40.8246
R6872 VSS.n4502 VSS.n1995 40.8246
R6873 VSS.n1990 VSS.n1963 40.8246
R6874 VSS.n1987 VSS.n1961 40.8246
R6875 VSS.n1986 VSS.n1985 40.8246
R6876 VSS.n1970 VSS.n1960 40.8246
R6877 VSS.n1972 VSS.n1967 40.8246
R6878 VSS.n1974 VSS.n1959 40.8246
R6879 VSS.n1976 VSS.n1968 40.8246
R6880 VSS.n1969 VSS.n1958 40.8246
R6881 VSS.n1983 VSS.n1982 40.8246
R6882 VSS.n1979 VSS.n1957 40.8246
R6883 VSS.n4526 VSS.n1953 40.8246
R6884 VSS.n1979 VSS.n1953 40.8246
R6885 VSS.n1982 VSS.n1957 40.8246
R6886 VSS.n1983 VSS.n1969 40.8246
R6887 VSS.n1976 VSS.n1958 40.8246
R6888 VSS.n1974 VSS.n1968 40.8246
R6889 VSS.n1972 VSS.n1959 40.8246
R6890 VSS.n1970 VSS.n1967 40.8246
R6891 VSS.n1985 VSS.n1960 40.8246
R6892 VSS.n1987 VSS.n1986 40.8246
R6893 VSS.n4008 VSS.n4007 40.8246
R6894 VSS.n2536 VSS.n1700 40.8246
R6895 VSS.n2538 VSS.n2537 40.8246
R6896 VSS.n2573 VSS.n1699 40.8246
R6897 VSS.n2572 VSS.n2571 40.8246
R6898 VSS.n2548 VSS.n1698 40.8246
R6899 VSS.n2550 VSS.n2549 40.8246
R6900 VSS.n2560 VSS.n1697 40.8246
R6901 VSS.n2559 VSS.n2558 40.8246
R6902 VSS.n3149 VSS.n1696 40.8246
R6903 VSS.n3148 VSS.n1703 40.8246
R6904 VSS.n3191 VSS.n3190 40.8246
R6905 VSS.n3372 VSS.n1694 40.8246
R6906 VSS.n3371 VSS.n3370 40.8246
R6907 VSS.n3245 VSS.n1693 40.8246
R6908 VSS.n3247 VSS.n3246 40.8246
R6909 VSS.n3254 VSS.n1692 40.8246
R6910 VSS.n3256 VSS.n3255 40.8246
R6911 VSS.n3263 VSS.n1691 40.8246
R6912 VSS.n3265 VSS.n3264 40.8246
R6913 VSS.n3381 VSS.n1690 40.8246
R6914 VSS.n3380 VSS.n1704 40.8246
R6915 VSS.n2394 VSS.n2393 40.8246
R6916 VSS.n2863 VSS.n1688 40.8246
R6917 VSS.n2865 VSS.n2864 40.8246
R6918 VSS.n2872 VSS.n1687 40.8246
R6919 VSS.n2874 VSS.n2873 40.8246
R6920 VSS.n2881 VSS.n1686 40.8246
R6921 VSS.n2883 VSS.n2882 40.8246
R6922 VSS.n2890 VSS.n1685 40.8246
R6923 VSS.n2892 VSS.n2891 40.8246
R6924 VSS.n2899 VSS.n1684 40.8246
R6925 VSS.n2898 VSS.n1705 40.8246
R6926 VSS.n2924 VSS.n2923 40.8246
R6927 VSS.n4625 VSS.n1682 40.8246
R6928 VSS.n4624 VSS.n4623 40.8246
R6929 VSS.n4404 VSS.n1681 40.8246
R6930 VSS.n4406 VSS.n4405 40.8246
R6931 VSS.n4413 VSS.n1680 40.8246
R6932 VSS.n4415 VSS.n4414 40.8246
R6933 VSS.n4422 VSS.n1679 40.8246
R6934 VSS.n4424 VSS.n4423 40.8246
R6935 VSS.n4431 VSS.n1678 40.8246
R6936 VSS.n4430 VSS.n1706 40.8246
R6937 VSS.n4689 VSS.n1670 40.8246
R6938 VSS.n4688 VSS.n1671 40.8246
R6939 VSS.n1783 VSS.n1782 40.8246
R6940 VSS.n1791 VSS.n1676 40.8246
R6941 VSS.n1796 VSS.n1784 40.8246
R6942 VSS.n1802 VSS.n1675 40.8246
R6943 VSS.n1807 VSS.n1785 40.8246
R6944 VSS.n1786 VSS.n1674 40.8246
R6945 VSS.n1825 VSS.n1824 40.8246
R6946 VSS.n1817 VSS.n1673 40.8246
R6947 VSS.n4686 VSS.n1707 40.8246
R6948 VSS.n2695 VSS.n2692 40.8246
R6949 VSS.n2696 VSS.n2695 40.8246
R6950 VSS.n2778 VSS.n2748 40.8246
R6951 VSS.n2750 VSS.n2748 40.8246
R6952 VSS.n3024 VSS.n2810 40.8246
R6953 VSS.n2812 VSS.n2810 40.8246
R6954 VSS.n4498 VSS.n1997 40.8246
R6955 VSS.n4499 VSS.n4498 40.8246
R6956 VSS.n4008 VSS.n1700 40.8246
R6957 VSS.n2538 VSS.n1699 40.8246
R6958 VSS.n2571 VSS.n1698 40.8246
R6959 VSS.n2550 VSS.n1697 40.8246
R6960 VSS.n2558 VSS.n1696 40.8246
R6961 VSS.n3191 VSS.n1694 40.8246
R6962 VSS.n3370 VSS.n1693 40.8246
R6963 VSS.n3247 VSS.n1692 40.8246
R6964 VSS.n3256 VSS.n1691 40.8246
R6965 VSS.n3265 VSS.n1690 40.8246
R6966 VSS.n2394 VSS.n1688 40.8246
R6967 VSS.n2865 VSS.n1687 40.8246
R6968 VSS.n2874 VSS.n1686 40.8246
R6969 VSS.n2883 VSS.n1685 40.8246
R6970 VSS.n2892 VSS.n1684 40.8246
R6971 VSS.n2924 VSS.n1682 40.8246
R6972 VSS.n4623 VSS.n1681 40.8246
R6973 VSS.n4406 VSS.n1680 40.8246
R6974 VSS.n4415 VSS.n1679 40.8246
R6975 VSS.n4424 VSS.n1678 40.8246
R6976 VSS.n4689 VSS.n4688 40.8246
R6977 VSS.n1782 VSS.n1676 40.8246
R6978 VSS.n1796 VSS.n1675 40.8246
R6979 VSS.n1807 VSS.n1674 40.8246
R6980 VSS.n1824 VSS.n1673 40.8246
R6981 VSS.n1817 VSS.n1707 40.8246
R6982 VSS.n1825 VSS.n1786 40.8246
R6983 VSS.n1802 VSS.n1785 40.8246
R6984 VSS.n1791 VSS.n1784 40.8246
R6985 VSS.n1783 VSS.n1671 40.8246
R6986 VSS.n1677 VSS.n1670 40.8246
R6987 VSS.n4431 VSS.n4430 40.8246
R6988 VSS.n4423 VSS.n4422 40.8246
R6989 VSS.n4414 VSS.n4413 40.8246
R6990 VSS.n4405 VSS.n4404 40.8246
R6991 VSS.n4625 VSS.n4624 40.8246
R6992 VSS.n2923 VSS.n1683 40.8246
R6993 VSS.n2899 VSS.n2898 40.8246
R6994 VSS.n2891 VSS.n2890 40.8246
R6995 VSS.n2882 VSS.n2881 40.8246
R6996 VSS.n2873 VSS.n2872 40.8246
R6997 VSS.n2864 VSS.n2863 40.8246
R6998 VSS.n2393 VSS.n1689 40.8246
R6999 VSS.n3381 VSS.n3380 40.8246
R7000 VSS.n3264 VSS.n3263 40.8246
R7001 VSS.n3255 VSS.n3254 40.8246
R7002 VSS.n3246 VSS.n3245 40.8246
R7003 VSS.n3372 VSS.n3371 40.8246
R7004 VSS.n3190 VSS.n1695 40.8246
R7005 VSS.n3149 VSS.n3148 40.8246
R7006 VSS.n2560 VSS.n2559 40.8246
R7007 VSS.n2549 VSS.n2548 40.8246
R7008 VSS.n2573 VSS.n2572 40.8246
R7009 VSS.n2537 VSS.n2536 40.8246
R7010 VSS.n4007 VSS.n1701 40.8246
R7011 VSS.n3187 VSS.n3155 40.8246
R7012 VSS.n3387 VSS.n2460 40.8246
R7013 VSS.n3388 VSS.n2460 40.8246
R7014 VSS.n2997 VSS.n2907 40.8246
R7015 VSS.n2999 VSS.n2929 40.8246
R7016 VSS.n1990 VSS.n1961 40.8246
R7017 VSS.n4524 VSS.n1963 40.8246
R7018 VSS.n1946 VSS.n1945 40.8246
R7019 VSS.n1942 VSS.n1893 40.8246
R7020 VSS.n1932 VSS.n1931 40.8246
R7021 VSS.n1928 VSS.n1906 40.8246
R7022 VSS.n1916 VSS.n1915 40.8246
R7023 VSS.n1918 VSS.n1917 40.8246
R7024 VSS.n1930 VSS.n1929 40.8246
R7025 VSS.n1904 VSS.n1903 40.8246
R7026 VSS.n1944 VSS.n1943 40.8246
R7027 VSS.n1948 VSS.n1947 40.8246
R7028 VSS.n2179 VSS.n158 40.8246
R7029 VSS.n3931 VSS.n658 40.8246
R7030 VSS.n2939 VSS.n672 40.8246
R7031 VSS.n4535 VSS.n864 40.8246
R7032 VSS.n5411 VSS.n5410 40.8246
R7033 VSS.n5407 VSS.n131 40.8246
R7034 VSS.n139 VSS.n138 40.8246
R7035 VSS.n5394 VSS.n140 40.8246
R7036 VSS.n155 VSS.n154 40.8246
R7037 VSS.n5118 VSS.n5117 40.8246
R7038 VSS.n5114 VSS.n631 40.8246
R7039 VSS.n639 VSS.n638 40.8246
R7040 VSS.n5101 VSS.n640 40.8246
R7041 VSS.n655 VSS.n654 40.8246
R7042 VSS.n2421 VSS.n2245 40.8246
R7043 VSS.n3906 VSS.n2246 40.8246
R7044 VSS.n3477 VSS.n3471 40.8246
R7045 VSS.n3488 VSS.n3487 40.8246
R7046 VSS.n3507 VSS.n3506 40.8246
R7047 VSS.n4890 VSS.n4889 40.8246
R7048 VSS.n4886 VSS.n838 40.8246
R7049 VSS.n846 VSS.n845 40.8246
R7050 VSS.n4873 VSS.n847 40.8246
R7051 VSS.n862 VSS.n861 40.8246
R7052 VSS.n4741 VSS.n1278 40.8246
R7053 VSS.n4768 VSS.n1279 40.8246
R7054 VSS.n1424 VSS.n1423 40.8246
R7055 VSS.n1429 VSS.n1428 40.8246
R7056 VSS.n1425 VSS.n1409 40.8246
R7057 VSS.n1483 VSS.n1482 40.8246
R7058 VSS.n1427 VSS.n1426 40.8246
R7059 VSS.n1431 VSS.n1430 40.8246
R7060 VSS.n1416 VSS.n1415 40.8246
R7061 VSS.n4770 VSS.n4769 40.8246
R7062 VSS.n4740 VSS.n4739 40.8246
R7063 VSS.n4862 VSS.n4861 40.8246
R7064 VSS.n860 VSS.n859 40.8246
R7065 VSS.n4875 VSS.n4874 40.8246
R7066 VSS.n844 VSS.n843 40.8246
R7067 VSS.n4888 VSS.n4887 40.8246
R7068 VSS.n4892 VSS.n4891 40.8246
R7069 VSS.n3509 VSS.n3508 40.8246
R7070 VSS.n3486 VSS.n3466 40.8246
R7071 VSS.n3485 VSS.n3484 40.8246
R7072 VSS.n3476 VSS.n3475 40.8246
R7073 VSS.n3908 VSS.n3907 40.8246
R7074 VSS.n2420 VSS.n663 40.8246
R7075 VSS.n5090 VSS.n5089 40.8246
R7076 VSS.n653 VSS.n652 40.8246
R7077 VSS.n5103 VSS.n5102 40.8246
R7078 VSS.n637 VSS.n636 40.8246
R7079 VSS.n5116 VSS.n5115 40.8246
R7080 VSS.n5120 VSS.n5119 40.8246
R7081 VSS.n5383 VSS.n5382 40.8246
R7082 VSS.n153 VSS.n152 40.8246
R7083 VSS.n5396 VSS.n5395 40.8246
R7084 VSS.n137 VSS.n136 40.8246
R7085 VSS.n5409 VSS.n5408 40.8246
R7086 VSS.n5413 VSS.n5412 40.8246
R7087 VSS.n5376 VSS.n157 40.8246
R7088 VSS.n5378 VSS.n161 40.8246
R7089 VSS.n5083 VSS.n657 40.8246
R7090 VSS.n5085 VSS.n661 40.8246
R7091 VSS.n5046 VSS.n671 40.8246
R7092 VSS.n5048 VSS.n674 40.8246
R7093 VSS.n4855 VSS.n863 40.8246
R7094 VSS.n4857 VSS.n867 40.8246
R7095 VSS.n1386 VSS.n1385 40.8246
R7096 VSS.n1558 VSS.n1557 40.8246
R7097 VSS.n5332 VSS.n243 40.8246
R7098 VSS.n5332 VSS.n242 40.8246
R7099 VSS.n3646 VSS.n3645 40.8246
R7100 VSS.n3647 VSS.n3646 40.8246
R7101 VSS.n5004 VSS.n5003 40.8246
R7102 VSS.n5004 VSS.n4977 40.8246
R7103 VSS.n1006 VSS.n272 40.8246
R7104 VSS.n1007 VSS.n1006 40.8246
R7105 VSS.n4316 VSS.n4230 39.8579
R7106 VSS.n4285 VSS.t72 39.0666
R7107 VSS.t73 VSS.t85 38.3621
R7108 VSS.n4784 VSS.n1245 37.6197
R7109 VSS.n5360 VSS.t32 36.9872
R7110 VSS.n4075 VSS.n69 36.9872
R7111 VSS.n5341 VSS.t32 36.9872
R7112 VSS.n4091 VSS.n27 36.9872
R7113 VSS.t35 VSS.n1672 36.9872
R7114 VSS.n4687 VSS.n1702 36.9872
R7115 VSS.n4258 VSS.n4254 36.563
R7116 VSS.n4257 VSS.n4254 36.563
R7117 VSS.n4277 VSS.n4276 36.563
R7118 VSS.n4277 VSS.n4237 36.563
R7119 VSS.n4075 VSS.n71 34.8534
R7120 VSS.n4091 VSS.n29 34.8534
R7121 VSS.n1826 VSS.n1702 34.8534
R7122 VSS.n4242 VSS.n4238 34.4123
R7123 VSS.n4256 VSS.n4238 34.4123
R7124 VSS.n4265 VSS.n4264 34.4123
R7125 VSS.n4264 VSS.t22 34.4123
R7126 VSS.n4263 VSS.n4262 34.4123
R7127 VSS.t22 VSS.n4263 34.4123
R7128 VSS.n4291 VSS.n4290 34.4123
R7129 VSS.n4292 VSS.n4291 34.4123
R7130 VSS.n4278 VSS.n4252 34.4123
R7131 VSS.t89 VSS.n4278 34.4123
R7132 VSS.n4280 VSS.n4279 34.4123
R7133 VSS.n4279 VSS.t89 34.4123
R7134 VSS.n5329 VSS.t32 33.3047
R7135 VSS.t74 VSS.t10 32.5716
R7136 VSS.n4857 VSS.n866 31.2084
R7137 VSS.n5378 VSS.n160 31.2084
R7138 VSS.n608 VSS.n183 31.2084
R7139 VSS.n194 VSS.n190 31.2084
R7140 VSS.n5343 VSS.n220 31.2084
R7141 VSS.n5006 VSS.n4968 31.2084
R7142 VSS.n5048 VSS.n669 31.2084
R7143 VSS.n5027 VSS.n697 31.2084
R7144 VSS.n994 VSS.n966 31.2084
R7145 VSS.n1033 VSS.n997 31.2084
R7146 VSS.n5334 VSS.n229 31.2084
R7147 VSS.n2207 VSS.n2206 31.2084
R7148 VSS.n3187 VSS.n2498 31.2084
R7149 VSS.n3419 VSS.n2463 31.2084
R7150 VSS.n3954 VSS.n2215 31.2084
R7151 VSS.n5085 VSS.n660 31.2084
R7152 VSS.n4560 VSS.n4527 31.2084
R7153 VSS.n2999 VSS.n2905 31.2084
R7154 VSS.n2964 VSS.n2963 31.2084
R7155 VSS.n4524 VSS.n1962 31.2084
R7156 VSS.n4315 VSS.n4314 30.8397
R7157 VSS.n1536 VSS.n1239 29.6284
R7158 VSS.n1485 VSS.n1227 29.6284
R7159 VSS.n4783 VSS.n4782 29.6284
R7160 VSS.n4783 VSS.n1248 29.6284
R7161 VSS.n1554 VSS.n1239 29.6284
R7162 VSS.n4306 VSS.n4305 28.3729
R7163 VSS.n4257 VSS.n4256 28.2149
R7164 VSS.t22 VSS.t11 25.3211
R7165 VSS.n5235 VSS.n270 24.3817
R7166 VSS.n5281 VSS.n271 24.3817
R7167 VSS.n5328 VSS.n5327 24.3817
R7168 VSS.n5330 VSS.n269 24.3817
R7169 VSS.t8 VSS.t26 23.8742
R7170 VSS.n4309 VSS.n4232 23.4005
R7171 VSS.n4303 VSS.n4232 23.4005
R7172 VSS.n4311 VSS.n4310 23.4005
R7173 VSS.n4312 VSS.n4311 23.4005
R7174 VSS.n4241 VSS.t14 21.5736
R7175 VSS.n4246 VSS.t18 21.5736
R7176 VSS.n4270 VSS.t24 21.5546
R7177 VSS.n4244 VSS.t17 21.4809
R7178 VSS.n4270 VSS.t13 21.4809
R7179 VSS.t32 VSS.n130 21.4062
R7180 VSS.n1844 VSS.t32 21.4062
R7181 VSS.n4298 VSS.n4297 18.1842
R7182 VSS.t38 VSS.t88 17.9811
R7183 VSS.n4191 VSS.n4173 17.4227
R7184 VSS.n5360 VSS.n69 16.36
R7185 VSS.n5341 VSS.n27 16.36
R7186 VSS.n4687 VSS.n1672 16.36
R7187 VSS.n1725 VSS.n1723 16.0005
R7188 VSS.n1723 VSS.n1720 16.0005
R7189 VSS.n1720 VSS.n1719 16.0005
R7190 VSS.n1719 VSS.n1716 16.0005
R7191 VSS.n1716 VSS.n1715 16.0005
R7192 VSS.n1715 VSS.n1712 16.0005
R7193 VSS.n1712 VSS.n1711 16.0005
R7194 VSS.n1711 VSS.n1253 16.0005
R7195 VSS.n2052 VSS.n2050 16.0005
R7196 VSS.n2050 VSS.n2047 16.0005
R7197 VSS.n2047 VSS.n2046 16.0005
R7198 VSS.n2046 VSS.n2043 16.0005
R7199 VSS.n2043 VSS.n2042 16.0005
R7200 VSS.n2042 VSS.n2039 16.0005
R7201 VSS.n2039 VSS.n2038 16.0005
R7202 VSS.n2038 VSS.n2035 16.0005
R7203 VSS.n2018 VSS.n2017 16.0005
R7204 VSS.n2017 VSS.n2014 16.0005
R7205 VSS.n2014 VSS.n2013 16.0005
R7206 VSS.n2013 VSS.n2010 16.0005
R7207 VSS.n2010 VSS.n2009 16.0005
R7208 VSS.n2009 VSS.n2006 16.0005
R7209 VSS.n2006 VSS.n1666 16.0005
R7210 VSS.n4709 VSS.n1666 16.0005
R7211 VSS.n4452 VSS.n4450 16.0005
R7212 VSS.n4450 VSS.n4447 16.0005
R7213 VSS.n4447 VSS.n4446 16.0005
R7214 VSS.n4446 VSS.n4443 16.0005
R7215 VSS.n4443 VSS.n4442 16.0005
R7216 VSS.n4442 VSS.n4439 16.0005
R7217 VSS.n4439 VSS.n4438 16.0005
R7218 VSS.n4438 VSS.n4435 16.0005
R7219 VSS.n2908 VSS.n1758 16.0005
R7220 VSS.n2911 VSS.n2908 16.0005
R7221 VSS.n2912 VSS.n2911 16.0005
R7222 VSS.n2915 VSS.n2912 16.0005
R7223 VSS.n2916 VSS.n2915 16.0005
R7224 VSS.n2919 VSS.n2916 16.0005
R7225 VSS.n2921 VSS.n2919 16.0005
R7226 VSS.n2922 VSS.n2921 16.0005
R7227 VSS.n2820 VSS.n2819 16.0005
R7228 VSS.n2823 VSS.n2820 16.0005
R7229 VSS.n2824 VSS.n2823 16.0005
R7230 VSS.n2827 VSS.n2824 16.0005
R7231 VSS.n2828 VSS.n2827 16.0005
R7232 VSS.n2831 VSS.n2828 16.0005
R7233 VSS.n2832 VSS.n2831 16.0005
R7234 VSS.n2835 VSS.n2832 16.0005
R7235 VSS.n2792 VSS.n2791 16.0005
R7236 VSS.n2791 VSS.n2788 16.0005
R7237 VSS.n2788 VSS.n2787 16.0005
R7238 VSS.n2787 VSS.n2784 16.0005
R7239 VSS.n2784 VSS.n2419 16.0005
R7240 VSS.n3426 VSS.n2419 16.0005
R7241 VSS.n3426 VSS.n3425 16.0005
R7242 VSS.n3425 VSS.n3424 16.0005
R7243 VSS.n2745 VSS.n2743 16.0005
R7244 VSS.n2743 VSS.n2740 16.0005
R7245 VSS.n2740 VSS.n2739 16.0005
R7246 VSS.n2739 VSS.n2736 16.0005
R7247 VSS.n2736 VSS.n2735 16.0005
R7248 VSS.n2735 VSS.n2732 16.0005
R7249 VSS.n2732 VSS.n2731 16.0005
R7250 VSS.n2731 VSS.n2464 16.0005
R7251 VSS.n2712 VSS.n2711 16.0005
R7252 VSS.n2711 VSS.n2708 16.0005
R7253 VSS.n2708 VSS.n2707 16.0005
R7254 VSS.n2707 VSS.n2704 16.0005
R7255 VSS.n2704 VSS.n2703 16.0005
R7256 VSS.n2703 VSS.n2700 16.0005
R7257 VSS.n2700 VSS.n2699 16.0005
R7258 VSS.n2699 VSS.n2493 16.0005
R7259 VSS.n2440 VSS.n2438 16.0005
R7260 VSS.n2438 VSS.n2435 16.0005
R7261 VSS.n2435 VSS.n2434 16.0005
R7262 VSS.n2434 VSS.n2431 16.0005
R7263 VSS.n2431 VSS.n2430 16.0005
R7264 VSS.n2430 VSS.n2427 16.0005
R7265 VSS.n2427 VSS.n2426 16.0005
R7266 VSS.n2426 VSS.n2424 16.0005
R7267 VSS.n2458 VSS.n2457 16.0005
R7268 VSS.n2457 VSS.n2454 16.0005
R7269 VSS.n2454 VSS.n2453 16.0005
R7270 VSS.n2453 VSS.n2450 16.0005
R7271 VSS.n2450 VSS.n2449 16.0005
R7272 VSS.n2449 VSS.n2446 16.0005
R7273 VSS.n2446 VSS.n2445 16.0005
R7274 VSS.n2445 VSS.n2442 16.0005
R7275 VSS.n2850 VSS.n2849 16.0005
R7276 VSS.n2849 VSS.n2846 16.0005
R7277 VSS.n2846 VSS.n2845 16.0005
R7278 VSS.n2845 VSS.n2842 16.0005
R7279 VSS.n2842 VSS.n2841 16.0005
R7280 VSS.n2841 VSS.n2838 16.0005
R7281 VSS.n2838 VSS.n2837 16.0005
R7282 VSS.n2837 VSS.n2322 16.0005
R7283 VSS.n3449 VSS.n3448 16.0005
R7284 VSS.n3452 VSS.n3449 16.0005
R7285 VSS.n3453 VSS.n3452 16.0005
R7286 VSS.n3456 VSS.n3453 16.0005
R7287 VSS.n3457 VSS.n3456 16.0005
R7288 VSS.n3460 VSS.n3457 16.0005
R7289 VSS.n3461 VSS.n3460 16.0005
R7290 VSS.n3464 VSS.n3461 16.0005
R7291 VSS.n4174 VSS.n126 16.0005
R7292 VSS.n4177 VSS.n4174 16.0005
R7293 VSS.n4178 VSS.n4177 16.0005
R7294 VSS.n4181 VSS.n4178 16.0005
R7295 VSS.n4182 VSS.n4181 16.0005
R7296 VSS.n4185 VSS.n4182 16.0005
R7297 VSS.n4186 VSS.n4185 16.0005
R7298 VSS.n4189 VSS.n4186 16.0005
R7299 VSS.n441 VSS.n440 16.0005
R7300 VSS.n444 VSS.n441 16.0005
R7301 VSS.n445 VSS.n444 16.0005
R7302 VSS.n448 VSS.n445 16.0005
R7303 VSS.n449 VSS.n448 16.0005
R7304 VSS.n452 VSS.n449 16.0005
R7305 VSS.n453 VSS.n452 16.0005
R7306 VSS.n456 VSS.n453 16.0005
R7307 VSS.n5481 VSS.n5480 16.0005
R7308 VSS.n5482 VSS.n5481 16.0005
R7309 VSS.n5482 VSS.n16 16.0005
R7310 VSS.n5488 VSS.n16 16.0005
R7311 VSS.n5489 VSS.n5488 16.0005
R7312 VSS.n5490 VSS.n5489 16.0005
R7313 VSS.n5490 VSS.n14 16.0005
R7314 VSS.n5496 VSS.n14 16.0005
R7315 VSS.n4173 VSS.n4172 16.0005
R7316 VSS.n4172 VSS.n4169 16.0005
R7317 VSS.n4169 VSS.n4168 16.0005
R7318 VSS.n4168 VSS.n4165 16.0005
R7319 VSS.n4165 VSS.n4164 16.0005
R7320 VSS.n4164 VSS.n4161 16.0005
R7321 VSS.n4161 VSS.n4160 16.0005
R7322 VSS.n4160 VSS.n4157 16.0005
R7323 VSS.n541 VSS.n540 16.0005
R7324 VSS.n540 VSS.n537 16.0005
R7325 VSS.n537 VSS.n536 16.0005
R7326 VSS.n536 VSS.n533 16.0005
R7327 VSS.n533 VSS.n532 16.0005
R7328 VSS.n532 VSS.n529 16.0005
R7329 VSS.n529 VSS.n528 16.0005
R7330 VSS.n528 VSS.n525 16.0005
R7331 VSS.n512 VSS.n457 16.0005
R7332 VSS.n512 VSS.n511 16.0005
R7333 VSS.n511 VSS.n510 16.0005
R7334 VSS.n510 VSS.n475 16.0005
R7335 VSS.n505 VSS.n475 16.0005
R7336 VSS.n505 VSS.n504 16.0005
R7337 VSS.n504 VSS.n503 16.0005
R7338 VSS.n503 VSS.n478 16.0005
R7339 VSS.n3725 VSS.n3711 16.0005
R7340 VSS.n3725 VSS.n3724 16.0005
R7341 VSS.n3724 VSS.n3723 16.0005
R7342 VSS.n3723 VSS.n3713 16.0005
R7343 VSS.n3718 VSS.n3713 16.0005
R7344 VSS.n3718 VSS.n3717 16.0005
R7345 VSS.n3717 VSS.n316 16.0005
R7346 VSS.n5229 VSS.n316 16.0005
R7347 VSS.n437 VSS.n436 16.0005
R7348 VSS.n436 VSS.n433 16.0005
R7349 VSS.n433 VSS.n432 16.0005
R7350 VSS.n432 VSS.n429 16.0005
R7351 VSS.n429 VSS.n428 16.0005
R7352 VSS.n428 VSS.n425 16.0005
R7353 VSS.n425 VSS.n424 16.0005
R7354 VSS.n424 VSS.n336 16.0005
R7355 VSS.n5177 VSS.n334 16.0005
R7356 VSS.n5183 VSS.n334 16.0005
R7357 VSS.n5184 VSS.n5183 16.0005
R7358 VSS.n5185 VSS.n5184 16.0005
R7359 VSS.n5185 VSS.n332 16.0005
R7360 VSS.n5191 VSS.n332 16.0005
R7361 VSS.n5192 VSS.n5191 16.0005
R7362 VSS.n5194 VSS.n5192 16.0005
R7363 VSS.n629 VSS.n628 16.0005
R7364 VSS.n628 VSS.n625 16.0005
R7365 VSS.n625 VSS.n624 16.0005
R7366 VSS.n624 VSS.n621 16.0005
R7367 VSS.n621 VSS.n620 16.0005
R7368 VSS.n620 VSS.n617 16.0005
R7369 VSS.n617 VSS.n616 16.0005
R7370 VSS.n616 VSS.n613 16.0005
R7371 VSS.n3734 VSS.n3733 16.0005
R7372 VSS.n3737 VSS.n3734 16.0005
R7373 VSS.n3738 VSS.n3737 16.0005
R7374 VSS.n3741 VSS.n3738 16.0005
R7375 VSS.n3742 VSS.n3741 16.0005
R7376 VSS.n3745 VSS.n3742 16.0005
R7377 VSS.n3746 VSS.n3745 16.0005
R7378 VSS.n3749 VSS.n3746 16.0005
R7379 VSS.n3785 VSS.n3782 16.0005
R7380 VSS.n3786 VSS.n3785 16.0005
R7381 VSS.n3789 VSS.n3786 16.0005
R7382 VSS.n3790 VSS.n3789 16.0005
R7383 VSS.n3793 VSS.n3790 16.0005
R7384 VSS.n3794 VSS.n3793 16.0005
R7385 VSS.n3797 VSS.n3794 16.0005
R7386 VSS.n3798 VSS.n3797 16.0005
R7387 VSS.n1187 VSS.n1186 16.0005
R7388 VSS.n1190 VSS.n1187 16.0005
R7389 VSS.n1191 VSS.n1190 16.0005
R7390 VSS.n1194 VSS.n1191 16.0005
R7391 VSS.n1195 VSS.n1194 16.0005
R7392 VSS.n1198 VSS.n1195 16.0005
R7393 VSS.n1200 VSS.n1198 16.0005
R7394 VSS.n1201 VSS.n1200 16.0005
R7395 VSS.n4760 VSS.n4759 16.0005
R7396 VSS.n4759 VSS.n4756 16.0005
R7397 VSS.n4756 VSS.n4755 16.0005
R7398 VSS.n4755 VSS.n4752 16.0005
R7399 VSS.n4752 VSS.n4751 16.0005
R7400 VSS.n4751 VSS.n4748 16.0005
R7401 VSS.n4748 VSS.n4747 16.0005
R7402 VSS.n4747 VSS.n4744 16.0005
R7403 VSS.n939 VSS.n938 16.0005
R7404 VSS.n942 VSS.n939 16.0005
R7405 VSS.n943 VSS.n942 16.0005
R7406 VSS.n946 VSS.n943 16.0005
R7407 VSS.n947 VSS.n946 16.0005
R7408 VSS.n950 VSS.n947 16.0005
R7409 VSS.n952 VSS.n950 16.0005
R7410 VSS.n953 VSS.n952 16.0005
R7411 VSS.n1580 VSS.n1577 16.0005
R7412 VSS.n1577 VSS.n1576 16.0005
R7413 VSS.n1576 VSS.n1573 16.0005
R7414 VSS.n1573 VSS.n1572 16.0005
R7415 VSS.n1572 VSS.n1569 16.0005
R7416 VSS.n1569 VSS.n1568 16.0005
R7417 VSS.n1568 VSS.n1565 16.0005
R7418 VSS.n1565 VSS.n1564 16.0005
R7419 VSS.n1340 VSS.n1338 16.0005
R7420 VSS.n1338 VSS.n1335 16.0005
R7421 VSS.n1335 VSS.n1334 16.0005
R7422 VSS.n1334 VSS.n1331 16.0005
R7423 VSS.n1331 VSS.n1330 16.0005
R7424 VSS.n1330 VSS.n1327 16.0005
R7425 VSS.n1327 VSS.n1326 16.0005
R7426 VSS.n1326 VSS.n1323 16.0005
R7427 VSS.n1102 VSS.n1037 16.0005
R7428 VSS.n1086 VSS.n1037 16.0005
R7429 VSS.n1095 VSS.n1086 16.0005
R7430 VSS.n1095 VSS.n1094 16.0005
R7431 VSS.n1094 VSS.n1093 16.0005
R7432 VSS.n1093 VSS.n1088 16.0005
R7433 VSS.n1088 VSS.n278 16.0005
R7434 VSS.n5321 VSS.n278 16.0005
R7435 VSS.n819 VSS.n818 16.0005
R7436 VSS.n818 VSS.n815 16.0005
R7437 VSS.n815 VSS.n814 16.0005
R7438 VSS.n814 VSS.n811 16.0005
R7439 VSS.n811 VSS.n810 16.0005
R7440 VSS.n810 VSS.n807 16.0005
R7441 VSS.n807 VSS.n725 16.0005
R7442 VSS.n4937 VSS.n725 16.0005
R7443 VSS.n4953 VSS.n4939 16.0005
R7444 VSS.n4953 VSS.n4952 16.0005
R7445 VSS.n4952 VSS.n4951 16.0005
R7446 VSS.n4951 VSS.n4941 16.0005
R7447 VSS.n4945 VSS.n4941 16.0005
R7448 VSS.n4945 VSS.n4944 16.0005
R7449 VSS.n4944 VSS.n292 16.0005
R7450 VSS.n5286 VSS.n292 16.0005
R7451 VSS.n837 VSS.n836 16.0005
R7452 VSS.n836 VSS.n833 16.0005
R7453 VSS.n833 VSS.n832 16.0005
R7454 VSS.n832 VSS.n829 16.0005
R7455 VSS.n829 VSS.n828 16.0005
R7456 VSS.n828 VSS.n825 16.0005
R7457 VSS.n825 VSS.n824 16.0005
R7458 VSS.n824 VSS.n821 16.0005
R7459 VSS.n1106 VSS.n1105 16.0005
R7460 VSS.n1109 VSS.n1106 16.0005
R7461 VSS.n1110 VSS.n1109 16.0005
R7462 VSS.n1113 VSS.n1110 16.0005
R7463 VSS.n1114 VSS.n1113 16.0005
R7464 VSS.n1117 VSS.n1114 16.0005
R7465 VSS.n1118 VSS.n1117 16.0005
R7466 VSS.n1121 VSS.n1118 16.0005
R7467 VSS.n1157 VSS.n1154 16.0005
R7468 VSS.n1158 VSS.n1157 16.0005
R7469 VSS.n1161 VSS.n1158 16.0005
R7470 VSS.n1162 VSS.n1161 16.0005
R7471 VSS.n1165 VSS.n1162 16.0005
R7472 VSS.n1166 VSS.n1165 16.0005
R7473 VSS.n1169 VSS.n1166 16.0005
R7474 VSS.n1172 VSS.n1169 16.0005
R7475 VSS.n3599 VSS.n3598 16.0005
R7476 VSS.n3598 VSS.n3583 16.0005
R7477 VSS.n3593 VSS.n3583 16.0005
R7478 VSS.n3593 VSS.n3592 16.0005
R7479 VSS.n3592 VSS.n3591 16.0005
R7480 VSS.n3591 VSS.n3586 16.0005
R7481 VSS.n3586 VSS.n297 16.0005
R7482 VSS.n5275 VSS.n297 16.0005
R7483 VSS.n3861 VSS.n2269 16.0005
R7484 VSS.n3861 VSS.n3860 16.0005
R7485 VSS.n3860 VSS.n3859 16.0005
R7486 VSS.n3859 VSS.n2271 16.0005
R7487 VSS.n3853 VSS.n2271 16.0005
R7488 VSS.n3853 VSS.n3852 16.0005
R7489 VSS.n3852 VSS.n3851 16.0005
R7490 VSS.n3851 VSS.n2273 16.0005
R7491 VSS.n3826 VSS.n3812 16.0005
R7492 VSS.n3826 VSS.n3825 16.0005
R7493 VSS.n3825 VSS.n3824 16.0005
R7494 VSS.n3824 VSS.n3814 16.0005
R7495 VSS.n3818 VSS.n3814 16.0005
R7496 VSS.n3818 VSS.n3817 16.0005
R7497 VSS.n3817 VSS.n311 16.0005
R7498 VSS.n5240 VSS.n311 16.0005
R7499 VSS.n3896 VSS.n2251 16.0005
R7500 VSS.n3896 VSS.n3895 16.0005
R7501 VSS.n3895 VSS.n3894 16.0005
R7502 VSS.n3894 VSS.n2253 16.0005
R7503 VSS.n3888 VSS.n2253 16.0005
R7504 VSS.n3888 VSS.n3887 16.0005
R7505 VSS.n3887 VSS.n3886 16.0005
R7506 VSS.n3886 VSS.n2255 16.0005
R7507 VSS.n3512 VSS.n2320 16.0005
R7508 VSS.n3518 VSS.n2320 16.0005
R7509 VSS.n3519 VSS.n3518 16.0005
R7510 VSS.n3520 VSS.n3519 16.0005
R7511 VSS.n3520 VSS.n2318 16.0005
R7512 VSS.n3525 VSS.n2318 16.0005
R7513 VSS.n3526 VSS.n3525 16.0005
R7514 VSS.n3526 VSS.n2308 16.0005
R7515 VSS.n3569 VSS.n3568 16.0005
R7516 VSS.n3569 VSS.n2306 16.0005
R7517 VSS.n3575 VSS.n2306 16.0005
R7518 VSS.n3576 VSS.n3575 16.0005
R7519 VSS.n3577 VSS.n3576 16.0005
R7520 VSS.n3577 VSS.n2304 16.0005
R7521 VSS.n3582 VSS.n2304 16.0005
R7522 VSS.n3601 VSS.n3582 16.0005
R7523 VSS.n5429 VSS.n125 16.0005
R7524 VSS.n5429 VSS.n5428 16.0005
R7525 VSS.n5428 VSS.n5427 16.0005
R7526 VSS.n5427 VSS.n5424 16.0005
R7527 VSS.n5424 VSS.n5423 16.0005
R7528 VSS.n5423 VSS.n5420 16.0005
R7529 VSS.n5420 VSS.n5419 16.0005
R7530 VSS.n5419 VSS.n5416 16.0005
R7531 VSS.n2105 VSS.n2081 16.0005
R7532 VSS.n2108 VSS.n2105 16.0005
R7533 VSS.n2109 VSS.n2108 16.0005
R7534 VSS.n2112 VSS.n2109 16.0005
R7535 VSS.n2113 VSS.n2112 16.0005
R7536 VSS.n4002 VSS.n2113 16.0005
R7537 VSS.n4002 VSS.n4001 16.0005
R7538 VSS.n4001 VSS.n4000 16.0005
R7539 VSS.n2514 VSS.n2513 16.0005
R7540 VSS.n2513 VSS.n2510 16.0005
R7541 VSS.n2510 VSS.n2509 16.0005
R7542 VSS.n2509 VSS.n2506 16.0005
R7543 VSS.n2506 VSS.n2505 16.0005
R7544 VSS.n2505 VSS.n2502 16.0005
R7545 VSS.n2502 VSS.n2501 16.0005
R7546 VSS.n2501 VSS.n2150 16.0005
R7547 VSS.n2168 VSS.n2166 16.0005
R7548 VSS.n2166 VSS.n2163 16.0005
R7549 VSS.n2163 VSS.n2162 16.0005
R7550 VSS.n2162 VSS.n2159 16.0005
R7551 VSS.n2159 VSS.n2158 16.0005
R7552 VSS.n2158 VSS.n2155 16.0005
R7553 VSS.n2155 VSS.n2154 16.0005
R7554 VSS.n2154 VSS.n2151 16.0005
R7555 VSS.n5136 VSS.n421 16.0005
R7556 VSS.n5136 VSS.n5135 16.0005
R7557 VSS.n5135 VSS.n5134 16.0005
R7558 VSS.n5134 VSS.n5131 16.0005
R7559 VSS.n5131 VSS.n5130 16.0005
R7560 VSS.n5130 VSS.n5127 16.0005
R7561 VSS.n5127 VSS.n5126 16.0005
R7562 VSS.n5126 VSS.n5123 16.0005
R7563 VSS.n3360 VSS.n3194 16.0005
R7564 VSS.n3360 VSS.n3359 16.0005
R7565 VSS.n3359 VSS.n3358 16.0005
R7566 VSS.n3358 VSS.n3196 16.0005
R7567 VSS.n3352 VSS.n3196 16.0005
R7568 VSS.n3352 VSS.n3351 16.0005
R7569 VSS.n3351 VSS.n3350 16.0005
R7570 VSS.n3350 VSS.n3198 16.0005
R7571 VSS.n3275 VSS.n2465 16.0005
R7572 VSS.n3276 VSS.n3275 16.0005
R7573 VSS.n3276 VSS.n3234 16.0005
R7574 VSS.n3282 VSS.n3234 16.0005
R7575 VSS.n3283 VSS.n3282 16.0005
R7576 VSS.n3284 VSS.n3283 16.0005
R7577 VSS.n3284 VSS.n3232 16.0005
R7578 VSS.n3289 VSS.n3232 16.0005
R7579 VSS.n3307 VSS.n3305 16.0005
R7580 VSS.n3305 VSS.n3302 16.0005
R7581 VSS.n3302 VSS.n3301 16.0005
R7582 VSS.n3301 VSS.n3298 16.0005
R7583 VSS.n3298 VSS.n3297 16.0005
R7584 VSS.n3297 VSS.n3294 16.0005
R7585 VSS.n3294 VSS.n3293 16.0005
R7586 VSS.n3293 VSS.n3290 16.0005
R7587 VSS.n4908 VSS.n806 16.0005
R7588 VSS.n4908 VSS.n4907 16.0005
R7589 VSS.n4907 VSS.n4906 16.0005
R7590 VSS.n4906 VSS.n4903 16.0005
R7591 VSS.n4903 VSS.n4902 16.0005
R7592 VSS.n4902 VSS.n4899 16.0005
R7593 VSS.n4899 VSS.n4898 16.0005
R7594 VSS.n4898 VSS.n4895 16.0005
R7595 VSS.n4613 VSS.n1831 16.0005
R7596 VSS.n4613 VSS.n4612 16.0005
R7597 VSS.n4612 VSS.n4611 16.0005
R7598 VSS.n4611 VSS.n1833 16.0005
R7599 VSS.n4605 VSS.n1833 16.0005
R7600 VSS.n4605 VSS.n4604 16.0005
R7601 VSS.n4604 VSS.n4603 16.0005
R7602 VSS.n4603 VSS.n1835 16.0005
R7603 VSS.n4389 VSS.n4367 16.0005
R7604 VSS.n4389 VSS.n4388 16.0005
R7605 VSS.n4388 VSS.n4387 16.0005
R7606 VSS.n4387 VSS.n4373 16.0005
R7607 VSS.n4382 VSS.n4373 16.0005
R7608 VSS.n4382 VSS.n4381 16.0005
R7609 VSS.n4381 VSS.n4380 16.0005
R7610 VSS.n4380 VSS.n4376 16.0005
R7611 VSS.n1885 VSS.n1883 16.0005
R7612 VSS.n1883 VSS.n1880 16.0005
R7613 VSS.n1880 VSS.n1879 16.0005
R7614 VSS.n1879 VSS.n1876 16.0005
R7615 VSS.n1876 VSS.n1875 16.0005
R7616 VSS.n1875 VSS.n1872 16.0005
R7617 VSS.n1872 VSS.n1871 16.0005
R7618 VSS.n1871 VSS.n1868 16.0005
R7619 VSS.n2658 VSS.n2656 16.0005
R7620 VSS.n2656 VSS.n2653 16.0005
R7621 VSS.n2653 VSS.n2652 16.0005
R7622 VSS.n2652 VSS.n2649 16.0005
R7623 VSS.n2649 VSS.n2648 16.0005
R7624 VSS.n2648 VSS.n2645 16.0005
R7625 VSS.n2645 VSS.n2644 16.0005
R7626 VSS.n2644 VSS.n2515 16.0005
R7627 VSS.n3128 VSS.n3127 16.0005
R7628 VSS.n3131 VSS.n3128 16.0005
R7629 VSS.n3132 VSS.n3131 16.0005
R7630 VSS.n3135 VSS.n3132 16.0005
R7631 VSS.n3136 VSS.n3135 16.0005
R7632 VSS.n3139 VSS.n3136 16.0005
R7633 VSS.n3140 VSS.n3139 16.0005
R7634 VSS.n3140 VSS.n2082 16.0005
R7635 VSS.n4707 VSS.n4704 16.0005
R7636 VSS.n4704 VSS.n4703 16.0005
R7637 VSS.n4703 VSS.n4700 16.0005
R7638 VSS.n4700 VSS.n4699 16.0005
R7639 VSS.n4699 VSS.n4696 16.0005
R7640 VSS.n4696 VSS.n4695 16.0005
R7641 VSS.n4695 VSS.n4692 16.0005
R7642 VSS.n4692 VSS.n4691 16.0005
R7643 VSS.n4723 VSS.n4722 16.0005
R7644 VSS.n4726 VSS.n4723 16.0005
R7645 VSS.n4727 VSS.n4726 16.0005
R7646 VSS.n4730 VSS.n4727 16.0005
R7647 VSS.n4731 VSS.n4730 16.0005
R7648 VSS.n4734 VSS.n4731 16.0005
R7649 VSS.n4736 VSS.n4734 16.0005
R7650 VSS.n4737 VSS.n4736 16.0005
R7651 VSS.n4777 VSS.n1255 16.0005
R7652 VSS.n1450 VSS.n1255 16.0005
R7653 VSS.n1453 VSS.n1450 16.0005
R7654 VSS.n1454 VSS.n1453 16.0005
R7655 VSS.n1457 VSS.n1454 16.0005
R7656 VSS.n1458 VSS.n1457 16.0005
R7657 VSS.n1461 VSS.n1458 16.0005
R7658 VSS.n1464 VSS.n1461 16.0005
R7659 VSS.n1479 VSS.n1476 16.0005
R7660 VSS.n1476 VSS.n1475 16.0005
R7661 VSS.n1475 VSS.n1472 16.0005
R7662 VSS.n1472 VSS.n1471 16.0005
R7663 VSS.n1471 VSS.n1468 16.0005
R7664 VSS.n1468 VSS.n1467 16.0005
R7665 VSS.n1467 VSS.n1321 16.0005
R7666 VSS.n1582 VSS.n1321 16.0005
R7667 VSS.n666 VSS.t32 15.1452
R7668 VSS.n2212 VSS.t32 15.1452
R7669 VSS.n5329 VSS.n6 14.7312
R7670 VSS.n4292 VSS.n4237 13.7528
R7671 VSS.n5480 VSS.n18 13.6894
R7672 VSS.n612 VSS.n437 13.6894
R7673 VSS.n5177 VSS.n5176 13.6894
R7674 VSS.n1186 VSS.n1183 13.6894
R7675 VSS.n938 VSS.n890 13.6894
R7676 VSS.n820 VSS.n819 13.6894
R7677 VSS.n4939 VSS.n4938 13.6894
R7678 VSS.n2269 VSS.n2268 13.6894
R7679 VSS.n3812 VSS.n3811 13.6894
R7680 VSS.n2018 VSS.n2005 13.5116
R7681 VSS.n4634 VSS.n1758 13.5116
R7682 VSS.n2792 VSS.n2779 13.5116
R7683 VSS.n3093 VSS.n2712 13.5116
R7684 VSS.n3127 VSS.n2583 13.5116
R7685 VSS.n2441 VSS.n2440 13.3338
R7686 VSS.n3422 VSS.n2458 13.3338
R7687 VSS.n5415 VSS.n126 13.3338
R7688 VSS.n5122 VSS.n629 13.3338
R7689 VSS.n4760 VSS.n4743 13.3338
R7690 VSS.n4894 VSS.n837 13.3338
R7691 VSS.n2423 VSS.n2251 13.3338
R7692 VSS.n3998 VSS.n125 13.3338
R7693 VSS.n4010 VSS.n2081 13.3338
R7694 VSS.n2169 VSS.n421 13.3338
R7695 VSS.n3194 VSS.n3193 13.3338
R7696 VSS.n2324 VSS.n806 13.3338
R7697 VSS.n2926 VSS.n1831 13.3338
R7698 VSS.n4708 VSS.n4707 13.3338
R7699 VSS.n4722 VSS.n1620 13.3338
R7700 VSS.n4271 VSS.n4241 12.1065
R7701 VSS.n1391 VSS.n1390 11.6369
R7702 VSS.n1394 VSS.n1391 11.6369
R7703 VSS.n1395 VSS.n1394 11.6369
R7704 VSS.n1398 VSS.n1395 11.6369
R7705 VSS.n1399 VSS.n1398 11.6369
R7706 VSS.n1402 VSS.n1399 11.6369
R7707 VSS.n1403 VSS.n1402 11.6369
R7708 VSS.n1406 VSS.n1403 11.6369
R7709 VSS.n4220 VSS.n4060 11.6369
R7710 VSS.n4214 VSS.n4060 11.6369
R7711 VSS.n4214 VSS.n4213 11.6369
R7712 VSS.n4213 VSS.n4212 11.6369
R7713 VSS.n4212 VSS.n4069 11.6369
R7714 VSS.n4206 VSS.n4069 11.6369
R7715 VSS.n4206 VSS.n4205 11.6369
R7716 VSS.n4205 VSS.n4204 11.6369
R7717 VSS.n4125 VSS.n4102 11.6369
R7718 VSS.n4125 VSS.n4124 11.6369
R7719 VSS.n4124 VSS.n4123 11.6369
R7720 VSS.n4123 VSS.n4103 11.6369
R7721 VSS.n4107 VSS.n4103 11.6369
R7722 VSS.n4115 VSS.n4107 11.6369
R7723 VSS.n4115 VSS.n4114 11.6369
R7724 VSS.n4114 VSS.n4113 11.6369
R7725 VSS.n4156 VSS.n4077 11.6369
R7726 VSS.n4150 VSS.n4077 11.6369
R7727 VSS.n4150 VSS.n4149 11.6369
R7728 VSS.n4149 VSS.n4148 11.6369
R7729 VSS.n4148 VSS.n4085 11.6369
R7730 VSS.n4142 VSS.n4085 11.6369
R7731 VSS.n4142 VSS.n4141 11.6369
R7732 VSS.n4141 VSS.n4140 11.6369
R7733 VSS.n4014 VSS.n2074 11.6369
R7734 VSS.n4021 VSS.n2074 11.6369
R7735 VSS.n4022 VSS.n4021 11.6369
R7736 VSS.n4023 VSS.n4022 11.6369
R7737 VSS.n4023 VSS.n2071 11.6369
R7738 VSS.n4029 VSS.n2071 11.6369
R7739 VSS.n4030 VSS.n4029 11.6369
R7740 VSS.n4032 VSS.n4030 11.6369
R7741 VSS.n4042 VSS.n2061 11.6369
R7742 VSS.n4049 VSS.n2061 11.6369
R7743 VSS.n4050 VSS.n4049 11.6369
R7744 VSS.n4051 VSS.n4050 11.6369
R7745 VSS.n4051 VSS.n2058 11.6369
R7746 VSS.n4058 VSS.n2058 11.6369
R7747 VSS.n4059 VSS.n4058 11.6369
R7748 VSS.n4222 VSS.n4059 11.6369
R7749 VSS.n2616 VSS.n2590 11.6369
R7750 VSS.n2616 VSS.n2615 11.6369
R7751 VSS.n2615 VSS.n2614 11.6369
R7752 VSS.n2614 VSS.n2594 11.6369
R7753 VSS.n2596 VSS.n2594 11.6369
R7754 VSS.n2605 VSS.n2596 11.6369
R7755 VSS.n2606 VSS.n2605 11.6369
R7756 VSS.n2606 VSS.n2078 11.6369
R7757 VSS.n4324 VSS.n4323 11.6369
R7758 VSS.n4325 VSS.n4324 11.6369
R7759 VSS.n4325 VSS.n1734 11.6369
R7760 VSS.n4640 VSS.n1734 11.6369
R7761 VSS.n4641 VSS.n4640 11.6369
R7762 VSS.n4642 VSS.n4641 11.6369
R7763 VSS.n4642 VSS.n1729 11.6369
R7764 VSS.n4650 VSS.n1729 11.6369
R7765 VSS.n4682 VSS.n4651 11.6369
R7766 VSS.n4676 VSS.n4651 11.6369
R7767 VSS.n4676 VSS.n4675 11.6369
R7768 VSS.n4675 VSS.n4674 11.6369
R7769 VSS.n4674 VSS.n4659 11.6369
R7770 VSS.n4668 VSS.n4659 11.6369
R7771 VSS.n4668 VSS.n4667 11.6369
R7772 VSS.n4667 VSS.n4666 11.6369
R7773 VSS.n1492 VSS.n1489 11.6369
R7774 VSS.n1493 VSS.n1492 11.6369
R7775 VSS.n1496 VSS.n1493 11.6369
R7776 VSS.n1497 VSS.n1496 11.6369
R7777 VSS.n1500 VSS.n1497 11.6369
R7778 VSS.n1501 VSS.n1500 11.6369
R7779 VSS.n1504 VSS.n1501 11.6369
R7780 VSS.n1505 VSS.n1504 11.6369
R7781 VSS.n1517 VSS.n1514 11.6369
R7782 VSS.n1518 VSS.n1517 11.6369
R7783 VSS.n1521 VSS.n1518 11.6369
R7784 VSS.n1522 VSS.n1521 11.6369
R7785 VSS.n1525 VSS.n1522 11.6369
R7786 VSS.n1526 VSS.n1525 11.6369
R7787 VSS.n1529 VSS.n1526 11.6369
R7788 VSS.n1530 VSS.n1529 11.6369
R7789 VSS.n1533 VSS.n1530 11.6369
R7790 VSS.n1551 VSS.n1548 11.6369
R7791 VSS.n1548 VSS.n1547 11.6369
R7792 VSS.n1547 VSS.n1544 11.6369
R7793 VSS.n1544 VSS.n1543 11.6369
R7794 VSS.n1543 VSS.n1540 11.6369
R7795 VSS.n1540 VSS.n1539 11.6369
R7796 VSS.n1539 VSS.n1220 11.6369
R7797 VSS.n4787 VSS.n1220 11.6369
R7798 VSS.n1552 VSS.n1551 11.0106
R7799 VSS.n1390 VSS.n1388 10.9261
R7800 VSS.n1534 VSS.n1533 10.9063
R7801 VSS.n4042 VSS.n4041 10.8998
R7802 VSS.t89 VSS.t7 10.8575
R7803 VSS.t12 VSS.t80 10.8575
R7804 VSS.n567 VSS.n541 10.3116
R7805 VSS.n524 VSS.n457 10.3116
R7806 VSS.n3711 VSS.n3630 10.3116
R7807 VSS.n3782 VSS.n3781 10.3116
R7808 VSS.n1581 VSS.n1580 10.3116
R7809 VSS.n1341 VSS.n1340 10.3116
R7810 VSS.n1173 VSS.n1102 10.3116
R7811 VSS.n1154 VSS.n1153 10.3116
R7812 VSS.n3600 VSS.n3599 10.3116
R7813 VSS.n3568 VSS.n3567 10.3116
R7814 VSS.n2053 VSS.n2052 10.1338
R7815 VSS.n4492 VSS.n4452 10.1338
R7816 VSS.n2819 VSS.n2809 10.1338
R7817 VSS.n2746 VSS.n2745 10.1338
R7818 VSS.n2659 VSS.n2658 10.1338
R7819 VSS.n4102 VSS.n4089 10.0853
R7820 VSS.n2623 VSS.n2590 10.0103
R7821 VSS.n4323 VSS.n4321 10.0103
R7822 VSS.n1726 VSS.n1725 9.95606
R7823 VSS.n2901 VSS.n2850 9.95606
R7824 VSS.n3448 VSS.n3446 9.95606
R7825 VSS.n440 VSS.n151 9.95606
R7826 VSS.n3733 VSS.n651 9.95606
R7827 VSS.n1105 VSS.n858 9.95606
R7828 VSS.n3512 VSS.n3511 9.95606
R7829 VSS.n3151 VSS.n2514 9.95606
R7830 VSS.n3966 VSS.n2168 9.95606
R7831 VSS.n3383 VSS.n2465 9.95606
R7832 VSS.n3308 VSS.n3307 9.95606
R7833 VSS.n4434 VSS.n4367 9.95606
R7834 VSS.n1886 VSS.n1885 9.95606
R7835 VSS.n4778 VSS.n4777 9.95606
R7836 VSS.n1480 VSS.n1479 9.95606
R7837 VSS.n4221 VSS.n4220 9.82676
R7838 VSS.n4014 VSS.n4013 9.82676
R7839 VSS.n4683 VSS.n4682 9.82676
R7840 VSS.n1489 VSS.n1488 9.82676
R7841 VSS.n1514 VSS.n1513 9.7416
R7842 VSS.n4273 VSS.n4272 9.29356
R7843 VSS.n4294 VSS.t5 8.7005
R7844 VSS.n4294 VSS.t29 8.7005
R7845 VSS.n4293 VSS.t3 8.7005
R7846 VSS.n4293 VSS.t1 8.7005
R7847 VSS.n4666 VSS.n1251 8.13406
R7848 VSS.n4032 VSS.n4031 8.00427
R7849 VSS.n4285 VSS.t19 7.95841
R7850 VSS.n1508 VSS.n1505 7.95163
R7851 VSS.n4778 VSS.n1253 7.11161
R7852 VSS.n3446 VSS.n2322 7.11161
R7853 VSS.n567 VSS.n456 7.11161
R7854 VSS.n525 VSS.n524 7.11161
R7855 VSS.n483 VSS.n478 7.11161
R7856 VSS.n5230 VSS.n5229 7.11161
R7857 VSS.n3781 VSS.n3749 7.11161
R7858 VSS.n3798 VSS.n3630 7.11161
R7859 VSS.n1564 VSS.n1341 7.11161
R7860 VSS.n1323 VSS.n1215 7.11161
R7861 VSS.n5322 VSS.n5321 7.11161
R7862 VSS.n1153 VSS.n1121 7.11161
R7863 VSS.n1173 VSS.n1172 7.11161
R7864 VSS.n5276 VSS.n5275 7.11161
R7865 VSS.n3567 VSS.n2308 7.11161
R7866 VSS.n3601 VSS.n3600 7.11161
R7867 VSS.n3966 VSS.n2150 7.11161
R7868 VSS.n3308 VSS.n3289 7.11161
R7869 VSS.n4376 VSS.n1886 7.11161
R7870 VSS.n1582 VSS.n1581 7.11161
R7871 VSS.n4272 VSS.n4271 7.102
R7872 VSS.n4781 VSS.n1251 7.06798
R7873 VSS.n1388 VSS.n1387 7.06798
R7874 VSS.n1535 VSS.n1534 6.94026
R7875 VSS.n1555 VSS.n1552 6.94026
R7876 VSS.n2035 VSS.n1726 6.93383
R7877 VSS.n4435 VSS.n4434 6.93383
R7878 VSS.n2901 VSS.n2835 6.93383
R7879 VSS.n3383 VSS.n2464 6.93383
R7880 VSS.n3511 VSS.n3464 6.93383
R7881 VSS.n2151 VSS.n151 6.93383
R7882 VSS.n3290 VSS.n651 6.93383
R7883 VSS.n1868 VSS.n858 6.93383
R7884 VSS.n3151 VSS.n2515 6.93383
R7885 VSS.n1480 VSS.n1464 6.93383
R7886 VSS.n4031 VSS.n2068 6.8987
R7887 VSS.n4041 VSS.n4040 6.8987
R7888 VSS.n1510 VSS.n1508 6.8987
R7889 VSS.n5051 VSS.n666 6.69939
R7890 VSS.n666 VSS.n129 6.69939
R7891 VSS.n3961 VSS.n2212 6.69939
R7892 VSS.n2212 VSS.n1841 6.69939
R7893 VSS.n1387 VSS.n1252 6.59682
R7894 VSS.n1556 VSS.n1555 6.47761
R7895 VSS.n4040 VSS.n2065 6.43882
R7896 VSS.n1513 VSS.n1383 6.43882
R7897 VSS.n1383 VSS.n1322 6.28553
R7898 VSS.n1537 VSS.n1381 6.16917
R7899 VSS.n1988 VSS.n1966 5.81868
R7900 VSS.n1971 VSS.n1966 5.81868
R7901 VSS.n1973 VSS.n1971 5.81868
R7902 VSS.n1975 VSS.n1973 5.81868
R7903 VSS.n1977 VSS.n1975 5.81868
R7904 VSS.n1978 VSS.n1977 5.81868
R7905 VSS.n1981 VSS.n1978 5.81868
R7906 VSS.n1981 VSS.n1980 5.81868
R7907 VSS.n5374 VSS.n5373 5.81868
R7908 VSS.n5373 VSS.n5371 5.81868
R7909 VSS.n5371 VSS.n169 5.81868
R7910 VSS.n173 VSS.n169 5.81868
R7911 VSS.n175 VSS.n173 5.81868
R7912 VSS.n177 VSS.n175 5.81868
R7913 VSS.n179 VSS.n177 5.81868
R7914 VSS.n5364 VSS.n179 5.81868
R7915 VSS.n4853 VSS.n4852 5.81868
R7916 VSS.n4852 VSS.n4850 5.81868
R7917 VSS.n4850 VSS.n875 5.81868
R7918 VSS.n879 VSS.n875 5.81868
R7919 VSS.n881 VSS.n879 5.81868
R7920 VSS.n883 VSS.n881 5.81868
R7921 VSS.n885 VSS.n883 5.81868
R7922 VSS.n4843 VSS.n885 5.81868
R7923 VSS.n992 VSS.n990 5.81868
R7924 VSS.n990 VSS.n968 5.81868
R7925 VSS.n973 VSS.n968 5.81868
R7926 VSS.n975 VSS.n973 5.81868
R7927 VSS.n977 VSS.n975 5.81868
R7928 VSS.n979 VSS.n977 5.81868
R7929 VSS.n980 VSS.n979 5.81868
R7930 VSS.n983 VSS.n980 5.81868
R7931 VSS.n983 VSS.n982 5.81868
R7932 VSS.n1026 VSS.n1000 5.81868
R7933 VSS.n1026 VSS.n1025 5.81868
R7934 VSS.n1025 VSS.n1002 5.81868
R7935 VSS.n1003 VSS.n1002 5.81868
R7936 VSS.n1017 VSS.n1003 5.81868
R7937 VSS.n1017 VSS.n1016 5.81868
R7938 VSS.n1016 VSS.n1005 5.81868
R7939 VSS.n1010 VSS.n1005 5.81868
R7940 VSS.n5044 VSS.n5043 5.81868
R7941 VSS.n5043 VSS.n5041 5.81868
R7942 VSS.n5041 VSS.n682 5.81868
R7943 VSS.n686 VSS.n682 5.81868
R7944 VSS.n688 VSS.n686 5.81868
R7945 VSS.n690 VSS.n688 5.81868
R7946 VSS.n692 VSS.n690 5.81868
R7947 VSS.n5034 VSS.n692 5.81868
R7948 VSS.n5023 VSS.n696 5.81868
R7949 VSS.n5023 VSS.n5022 5.81868
R7950 VSS.n5022 VSS.n5020 5.81868
R7951 VSS.n5020 VSS.n707 5.81868
R7952 VSS.n711 VSS.n707 5.81868
R7953 VSS.n713 VSS.n711 5.81868
R7954 VSS.n715 VSS.n713 5.81868
R7955 VSS.n717 VSS.n715 5.81868
R7956 VSS.n5013 VSS.n717 5.81868
R7957 VSS.n5081 VSS.n5080 5.81868
R7958 VSS.n5080 VSS.n5078 5.81868
R7959 VSS.n5078 VSS.n5060 5.81868
R7960 VSS.n5064 VSS.n5060 5.81868
R7961 VSS.n5066 VSS.n5064 5.81868
R7962 VSS.n5068 VSS.n5066 5.81868
R7963 VSS.n5070 VSS.n5068 5.81868
R7964 VSS.n5071 VSS.n5070 5.81868
R7965 VSS.n5353 VSS.n195 5.81868
R7966 VSS.n208 VSS.n195 5.81868
R7967 VSS.n210 VSS.n208 5.81868
R7968 VSS.n212 VSS.n210 5.81868
R7969 VSS.n213 VSS.n212 5.81868
R7970 VSS.n215 VSS.n213 5.81868
R7971 VSS.n215 VSS.n214 5.81868
R7972 VSS.n214 VSS.n203 5.81868
R7973 VSS.n5346 VSS.n203 5.81868
R7974 VSS.n3663 VSS.n3632 5.81868
R7975 VSS.n3663 VSS.n3662 5.81868
R7976 VSS.n3662 VSS.n3638 5.81868
R7977 VSS.n3639 VSS.n3638 5.81868
R7978 VSS.n3654 VSS.n3639 5.81868
R7979 VSS.n3654 VSS.n3653 5.81868
R7980 VSS.n3653 VSS.n3641 5.81868
R7981 VSS.n3642 VSS.n3641 5.81868
R7982 VSS.n4992 VSS.n4983 5.81868
R7983 VSS.n4992 VSS.n4991 5.81868
R7984 VSS.n4991 VSS.n4989 5.81868
R7985 VSS.n4989 VSS.n4987 5.81868
R7986 VSS.n4987 VSS.n4985 5.81868
R7987 VSS.n4985 VSS.n4978 5.81868
R7988 VSS.n4998 VSS.n4978 5.81868
R7989 VSS.n5000 VSS.n4998 5.81868
R7990 VSS.n258 VSS.n249 5.81868
R7991 VSS.n258 VSS.n257 5.81868
R7992 VSS.n257 VSS.n255 5.81868
R7993 VSS.n255 VSS.n253 5.81868
R7994 VSS.n253 VSS.n251 5.81868
R7995 VSS.n251 VSS.n244 5.81868
R7996 VSS.n264 VSS.n244 5.81868
R7997 VSS.n266 VSS.n264 5.81868
R7998 VSS.n604 VSS.n573 5.81868
R7999 VSS.n604 VSS.n603 5.81868
R8000 VSS.n603 VSS.n601 5.81868
R8001 VSS.n601 VSS.n583 5.81868
R8002 VSS.n587 VSS.n583 5.81868
R8003 VSS.n589 VSS.n587 5.81868
R8004 VSS.n591 VSS.n589 5.81868
R8005 VSS.n593 VSS.n591 5.81868
R8006 VSS.n594 VSS.n593 5.81868
R8007 VSS.n3183 VSS.n3182 5.81868
R8008 VSS.n3182 VSS.n3181 5.81868
R8009 VSS.n3181 VSS.n3158 5.81868
R8010 VSS.n3160 VSS.n3158 5.81868
R8011 VSS.n3163 VSS.n3160 5.81868
R8012 VSS.n3171 VSS.n3163 5.81868
R8013 VSS.n3171 VSS.n3170 5.81868
R8014 VSS.n3170 VSS.n3169 5.81868
R8015 VSS.n2194 VSS.n2187 5.81868
R8016 VSS.n2194 VSS.n2193 5.81868
R8017 VSS.n2193 VSS.n2191 5.81868
R8018 VSS.n2191 VSS.n2189 5.81868
R8019 VSS.n2189 VSS.n2180 5.81868
R8020 VSS.n2200 VSS.n2180 5.81868
R8021 VSS.n2201 VSS.n2200 5.81868
R8022 VSS.n2202 VSS.n2201 5.81868
R8023 VSS.n3401 VSS.n3399 5.81868
R8024 VSS.n3403 VSS.n3401 5.81868
R8025 VSS.n3405 VSS.n3403 5.81868
R8026 VSS.n3407 VSS.n3405 5.81868
R8027 VSS.n3409 VSS.n3407 5.81868
R8028 VSS.n3410 VSS.n3409 5.81868
R8029 VSS.n3412 VSS.n3410 5.81868
R8030 VSS.n3412 VSS.n3411 5.81868
R8031 VSS.n3947 VSS.n3924 5.81868
R8032 VSS.n3947 VSS.n3946 5.81868
R8033 VSS.n3946 VSS.n3926 5.81868
R8034 VSS.n3927 VSS.n3926 5.81868
R8035 VSS.n3938 VSS.n3927 5.81868
R8036 VSS.n3938 VSS.n3937 5.81868
R8037 VSS.n3937 VSS.n3929 5.81868
R8038 VSS.n3930 VSS.n3929 5.81868
R8039 VSS.n4548 VSS.n4541 5.81868
R8040 VSS.n4548 VSS.n4547 5.81868
R8041 VSS.n4547 VSS.n4545 5.81868
R8042 VSS.n4545 VSS.n4543 5.81868
R8043 VSS.n4543 VSS.n4536 5.81868
R8044 VSS.n4554 VSS.n4536 5.81868
R8045 VSS.n4555 VSS.n4554 5.81868
R8046 VSS.n4556 VSS.n4555 5.81868
R8047 VSS.n2995 VSS.n2994 5.81868
R8048 VSS.n2994 VSS.n2992 5.81868
R8049 VSS.n2992 VSS.n2972 5.81868
R8050 VSS.n2976 VSS.n2972 5.81868
R8051 VSS.n2978 VSS.n2976 5.81868
R8052 VSS.n2980 VSS.n2978 5.81868
R8053 VSS.n2982 VSS.n2980 5.81868
R8054 VSS.n2985 VSS.n2982 5.81868
R8055 VSS.n2959 VSS.n2933 5.81868
R8056 VSS.n2934 VSS.n2933 5.81868
R8057 VSS.n2951 VSS.n2934 5.81868
R8058 VSS.n2951 VSS.n2950 5.81868
R8059 VSS.n2950 VSS.n2936 5.81868
R8060 VSS.n2937 VSS.n2936 5.81868
R8061 VSS.n2942 VSS.n2937 5.81868
R8062 VSS.n2942 VSS.n2941 5.81868
R8063 VSS.n4503 VSS.n1996 5.81868
R8064 VSS.n4504 VSS.n4503 5.81868
R8065 VSS.n4504 VSS.n1994 5.81868
R8066 VSS.n4510 VSS.n1994 5.81868
R8067 VSS.n4511 VSS.n4510 5.81868
R8068 VSS.n4511 VSS.n1992 5.81868
R8069 VSS.n4517 VSS.n1992 5.81868
R8070 VSS.n4518 VSS.n4517 5.81868
R8071 VSS.n2776 VSS.n2749 5.81868
R8072 VSS.n2770 VSS.n2749 5.81868
R8073 VSS.n2770 VSS.n2769 5.81868
R8074 VSS.n2769 VSS.n2752 5.81868
R8075 VSS.n2753 VSS.n2752 5.81868
R8076 VSS.n2761 VSS.n2753 5.81868
R8077 VSS.n2761 VSS.n2760 5.81868
R8078 VSS.n2760 VSS.n2755 5.81868
R8079 VSS.n3022 VSS.n2811 5.81868
R8080 VSS.n3016 VSS.n2811 5.81868
R8081 VSS.n3016 VSS.n3015 5.81868
R8082 VSS.n3015 VSS.n2814 5.81868
R8083 VSS.n2815 VSS.n2814 5.81868
R8084 VSS.n3007 VSS.n2815 5.81868
R8085 VSS.n3007 VSS.n3006 5.81868
R8086 VSS.n3006 VSS.n2817 5.81868
R8087 VSS.n2687 VSS.n2669 5.81868
R8088 VSS.n2687 VSS.n2686 5.81868
R8089 VSS.n2686 VSS.n2685 5.81868
R8090 VSS.n2685 VSS.n2670 5.81868
R8091 VSS.n2672 VSS.n2670 5.81868
R8092 VSS.n2675 VSS.n2672 5.81868
R8093 VSS.n2677 VSS.n2675 5.81868
R8094 VSS.n2677 VSS.n2676 5.81868
R8095 VSS.n1000 VSS.n956 5.51409
R8096 VSS.n3669 VSS.n3632 5.51409
R8097 VSS.n4983 VSS.n4967 5.51409
R8098 VSS.n249 VSS.n233 5.51409
R8099 VSS.n493 VSS.n492 5.50178
R8100 VSS.n3644 VSS.n313 5.50178
R8101 VSS.n5002 VSS.n294 5.50178
R8102 VSS.n1008 VSS.n275 5.50178
R8103 VSS.n4789 VSS.n4788 5.50178
R8104 VSS.n2694 VSS.n2693 5.47847
R8105 VSS.n3062 VSS.n3061 5.47847
R8106 VSS.n3027 VSS.n3026 5.47847
R8107 VSS.n4493 VSS.n1998 5.47847
R8108 VSS.n4321 VSS.n4320 5.47847
R8109 VSS.n982 VSS.n959 5.46332
R8110 VSS.n5013 VSS.n5012 5.46332
R8111 VSS.n5346 VSS.n5345 5.46332
R8112 VSS.n594 VSS.n230 5.46332
R8113 VSS.n2187 VSS.n2186 5.46332
R8114 VSS.n3924 VSS.n3921 5.46332
R8115 VSS.n4541 VSS.n1951 5.46332
R8116 VSS.n2960 VSS.n2959 5.46332
R8117 VSS.n5498 VSS.n13 5.22944
R8118 VSS.n5331 VSS.n268 5.22944
R8119 VSS.n5238 VSS.n312 5.22944
R8120 VSS.n5284 VSS.n293 5.22944
R8121 VSS.n1202 VSS.n273 5.22944
R8122 VSS.n2624 VSS.n2623 5.20728
R8123 VSS.n3094 VSS.n2697 5.20728
R8124 VSS.n3059 VSS.n3058 5.20728
R8125 VSS.n4635 VSS.n1757 5.20728
R8126 VSS.n4497 VSS.n2000 5.20728
R8127 VSS.n1999 VSS.n1996 4.97828
R8128 VSS.n2777 VSS.n2776 4.97828
R8129 VSS.n3023 VSS.n3022 4.97828
R8130 VSS.n2669 VSS.n2665 4.97828
R8131 VSS.n4288 VSS.n4287 4.95702
R8132 VSS.n1989 VSS.n1988 4.91363
R8133 VSS.n5374 VSS.n159 4.91363
R8134 VSS.n4853 VSS.n865 4.91363
R8135 VSS.n5044 VSS.n673 4.91363
R8136 VSS.n5081 VSS.n659 4.91363
R8137 VSS.n3183 VSS.n2494 4.91363
R8138 VSS.n3399 VSS.n2459 4.91363
R8139 VSS.n2995 VSS.n2906 4.91363
R8140 VSS.n993 VSS.n992 4.90491
R8141 VSS.n5028 VSS.n696 4.90491
R8142 VSS.n5354 VSS.n5353 4.90491
R8143 VSS.n609 VSS.n573 4.90491
R8144 VSS.n4307 VSS.n4235 4.71144
R8145 VSS.n4247 VSS 4.42669
R8146 VSS.n4780 VSS.n4779 4.24099
R8147 VSS.n2115 VSS.n2114 4.13942
R8148 VSS.n1980 VSS.n1955 4.06728
R8149 VSS.n3169 VSS.n3168 4.06728
R8150 VSS.n3411 VSS.n2216 4.06728
R8151 VSS.n2985 VSS.n2984 4.06728
R8152 VSS.n5364 VSS.n5363 4.0419
R8153 VSS.n4843 VSS.n4842 4.0419
R8154 VSS.n5034 VSS.n5033 4.0419
R8155 VSS.n5071 VSS.n191 4.0419
R8156 VSS.n11 VSS.n10 4.03114
R8157 VSS.n5505 VSS.n5504 4.03114
R8158 VSS.n5509 VSS.n8 4.03114
R8159 VSS.n5510 VSS.n4 4.03114
R8160 VSS.n5515 VSS.n5514 4.03114
R8161 VSS.n486 VSS.n1 4.03114
R8162 VSS.n488 VSS.n487 4.03114
R8163 VSS.n498 VSS.n482 4.03114
R8164 VSS.n5198 VSS.n330 4.03114
R8165 VSS.n5200 VSS.n5199 4.03114
R8166 VSS.n5207 VSS.n326 4.03114
R8167 VSS.n5206 VSS.n324 4.03114
R8168 VSS.n5213 VSS.n323 4.03114
R8169 VSS.n5222 VSS.n321 4.03114
R8170 VSS.n5221 VSS.n319 4.03114
R8171 VSS.n318 VSS.n315 4.03114
R8172 VSS.n5244 VSS.n309 4.03114
R8173 VSS.n5246 VSS.n5245 4.03114
R8174 VSS.n5253 VSS.n307 4.03114
R8175 VSS.n5252 VSS.n305 4.03114
R8176 VSS.n5259 VSS.n304 4.03114
R8177 VSS.n5268 VSS.n302 4.03114
R8178 VSS.n5267 VSS.n300 4.03114
R8179 VSS.n299 VSS.n296 4.03114
R8180 VSS.n5290 VSS.n290 4.03114
R8181 VSS.n5292 VSS.n5291 4.03114
R8182 VSS.n5299 VSS.n288 4.03114
R8183 VSS.n5298 VSS.n286 4.03114
R8184 VSS.n5305 VSS.n285 4.03114
R8185 VSS.n5314 VSS.n283 4.03114
R8186 VSS.n5313 VSS.n281 4.03114
R8187 VSS.n280 VSS.n277 4.03114
R8188 VSS.n4819 VSS.n1204 4.03114
R8189 VSS.n4818 VSS.n1205 4.03114
R8190 VSS.n4814 VSS.n4813 4.03114
R8191 VSS.n4811 VSS.n4810 4.03114
R8192 VSS.n4807 VSS.n1209 4.03114
R8193 VSS.n4802 VSS.n4801 4.03114
R8194 VSS.n4798 VSS.n4797 4.03114
R8195 VSS.n4794 VSS.n1214 4.03114
R8196 VSS VSS.n5519 3.97667
R8197 VSS VSS.n5214 3.97667
R8198 VSS VSS.n5260 3.97667
R8199 VSS VSS.n5306 3.97667
R8200 VSS.n1213 VSS 3.97667
R8201 VSS.n2442 VSS.n2441 3.73383
R8202 VSS.n4190 VSS.n4189 3.73383
R8203 VSS.n5497 VSS.n5496 3.73383
R8204 VSS.n4157 VSS.n18 3.73383
R8205 VSS.n5176 VSS.n336 3.73383
R8206 VSS.n5194 VSS.n5193 3.73383
R8207 VSS.n613 VSS.n612 3.73383
R8208 VSS.n1203 VSS.n1201 3.73383
R8209 VSS.n4744 VSS.n890 3.73383
R8210 VSS.n1183 VSS.n953 3.73383
R8211 VSS.n4938 VSS.n4937 3.73383
R8212 VSS.n5286 VSS.n5285 3.73383
R8213 VSS.n821 VSS.n820 3.73383
R8214 VSS.n3811 VSS.n2273 3.73383
R8215 VSS.n5240 VSS.n5239 3.73383
R8216 VSS.n2268 VSS.n2255 3.73383
R8217 VSS.n4000 VSS.n3998 3.73383
R8218 VSS.n3198 VSS.n2169 3.73383
R8219 VSS.n2324 VSS.n1835 3.73383
R8220 VSS.n4691 VSS.n1620 3.73383
R8221 VSS.n4779 VSS.n1252 3.6913
R8222 VSS.t75 VSS.t16 3.61773
R8223 VSS.n2115 VSS.n2065 3.6029
R8224 VSS.n4709 VSS.n4708 3.55606
R8225 VSS.n2926 VSS.n2922 3.55606
R8226 VSS.n3424 VSS.n3422 3.55606
R8227 VSS.n3193 VSS.n2493 3.55606
R8228 VSS.n2424 VSS.n2423 3.55606
R8229 VSS.n5416 VSS.n5415 3.55606
R8230 VSS.n5123 VSS.n5122 3.55606
R8231 VSS.n4895 VSS.n4894 3.55606
R8232 VSS.n4010 VSS.n2082 3.55606
R8233 VSS.n4743 VSS.n4737 3.55606
R8234 VSS.n4842 VSS.n4841 3.53424
R8235 VSS.n959 VSS.n958 3.53424
R8236 VSS.n1034 VSS.n956 3.53424
R8237 VSS.n5033 VSS.n5032 3.53424
R8238 VSS.n5358 VSS.n191 3.53424
R8239 VSS.n5345 VSS.n219 3.53424
R8240 VSS.n3670 VSS.n3669 3.53424
R8241 VSS.n5012 VSS.n5011 3.53424
R8242 VSS.n5007 VSS.n4967 3.53424
R8243 VSS.n5339 VSS.n230 3.53424
R8244 VSS.n5335 VSS.n233 3.53424
R8245 VSS.n5363 VSS.n5362 3.53424
R8246 VSS.n3168 VSS.n2208 3.53424
R8247 VSS.n2186 VSS.n2172 3.53424
R8248 VSS.n3959 VSS.n2216 3.53424
R8249 VSS.n3955 VSS.n3921 3.53424
R8250 VSS.n1955 VSS.n1954 3.53424
R8251 VSS.n4561 VSS.n1951 3.53424
R8252 VSS.n2984 VSS.n2983 3.53424
R8253 VSS.n2960 VSS.n2330 3.53424
R8254 VSS.n993 VSS.n888 3.29866
R8255 VSS.n1178 VSS.n1034 3.29866
R8256 VSS.n5029 VSS.n5028 3.29866
R8257 VSS.n5355 VSS.n5354 3.29866
R8258 VSS.n3806 VSS.n3670 3.29866
R8259 VSS.n5008 VSS.n5007 3.29866
R8260 VSS.n5336 VSS.n5335 3.29866
R8261 VSS.n610 VSS.n609 3.29866
R8262 VSS.n3964 VSS.n2172 3.29866
R8263 VSS.n3956 VSS.n3955 3.29866
R8264 VSS.n4562 VSS.n4561 3.29866
R8265 VSS.n3444 VSS.n2330 3.29866
R8266 VSS.n4229 VSS.n4228 3.22364
R8267 VSS.n888 VSS.n887 3.22013
R8268 VSS.n5029 VSS.n694 3.22013
R8269 VSS.n5355 VSS.n192 3.22013
R8270 VSS.n611 VSS.n610 3.22013
R8271 VSS.n4274 VSS.n4273 3.15497
R8272 VSS.n955 VSS.n954 3.1416
R8273 VSS.n3807 VSS.n3631 3.1416
R8274 VSS.n5010 VSS.n719 3.1416
R8275 VSS.n5338 VSS.n231 3.1416
R8276 VSS.n4275 VSS.n4236 3.1005
R8277 VSS.n4308 VSS.n4307 2.86813
R8278 VSS.n5498 VSS.n5497 2.83284
R8279 VSS.n5193 VSS.n268 2.83284
R8280 VSS.n5239 VSS.n5238 2.83284
R8281 VSS.n5285 VSS.n5284 2.83284
R8282 VSS.n1203 VSS.n1202 2.83284
R8283 VSS.n4315 VSS.n4231 2.82934
R8284 VSS.n2624 VSS.n2583 2.82084
R8285 VSS.n3094 VSS.n3093 2.82084
R8286 VSS.n3058 VSS.n2779 2.82084
R8287 VSS.n4635 VSS.n4634 2.82084
R8288 VSS.n2005 VSS.n2000 2.82084
R8289 VSS.n5331 VSS.n267 2.77837
R8290 VSS.n3643 VSS.n312 2.77837
R8291 VSS.n5001 VSS.n293 2.77837
R8292 VSS.n1009 VSS.n273 2.77837
R8293 VSS.n2697 VSS.n2665 2.7666
R8294 VSS.n3059 VSS.n2777 2.7666
R8295 VSS.n3023 VSS.n1757 2.7666
R8296 VSS.n4497 VSS.n1999 2.7666
R8297 VSS.n3154 VSS.n3152 2.73369
R8298 VSS.n3386 VSS.n3384 2.73369
R8299 VSS.n2903 VSS.n2902 2.73369
R8300 VSS.n4433 VSS.n1965 2.73369
R8301 VSS.n4685 VSS.n4684 2.73369
R8302 VSS.n5380 VSS.n5379 2.73369
R8303 VSS.n5087 VSS.n5086 2.73369
R8304 VSS.n5049 VSS.n670 2.73369
R8305 VSS.n4859 VSS.n4858 2.73369
R8306 VSS.n1487 VSS.n1407 2.73369
R8307 VSS.n492 VSS.n267 2.7239
R8308 VSS.n3644 VSS.n3643 2.7239
R8309 VSS.n5002 VSS.n5001 2.7239
R8310 VSS.n1009 VSS.n1008 2.7239
R8311 VSS.n3124 VSS.n3123 2.71236
R8312 VSS.n2630 VSS.n2585 2.71236
R8313 VSS.n3117 VSS.n2633 2.71236
R8314 VSS.n3116 VSS.n2634 2.71236
R8315 VSS.n3113 VSS.n3112 2.71236
R8316 VSS.n2639 VSS.n2635 2.71236
R8317 VSS.n3106 VSS.n2642 2.71236
R8318 VSS.n3105 VSS.n3103 2.71236
R8319 VSS.n3102 VSS.n3101 2.71236
R8320 VSS.n2694 VSS.n2665 2.71236
R8321 VSS.n3091 VSS.n3088 2.71236
R8322 VSS.n2717 VSS.n2713 2.71236
R8323 VSS.n3082 VSS.n2720 2.71236
R8324 VSS.n3081 VSS.n2721 2.71236
R8325 VSS.n3078 VSS.n3077 2.71236
R8326 VSS.n2726 VSS.n2722 2.71236
R8327 VSS.n3071 VSS.n2729 2.71236
R8328 VSS.n3070 VSS.n3068 2.71236
R8329 VSS.n3067 VSS.n3066 2.71236
R8330 VSS.n3061 VSS.n2777 2.71236
R8331 VSS.n2796 VSS.n2795 2.71236
R8332 VSS.n3051 VSS.n2797 2.71236
R8333 VSS.n3050 VSS.n3047 2.71236
R8334 VSS.n3046 VSS.n2798 2.71236
R8335 VSS.n3043 VSS.n3042 2.71236
R8336 VSS.n2805 VSS.n2799 2.71236
R8337 VSS.n3036 VSS.n2808 2.71236
R8338 VSS.n3035 VSS.n3033 2.71236
R8339 VSS.n3032 VSS.n3031 2.71236
R8340 VSS.n3026 VSS.n3023 2.71236
R8341 VSS.n4632 VSS.n1759 2.71236
R8342 VSS.n4462 VSS.n4461 2.71236
R8343 VSS.n4471 VSS.n4460 2.71236
R8344 VSS.n4472 VSS.n4458 2.71236
R8345 VSS.n4476 VSS.n4475 2.71236
R8346 VSS.n4482 VSS.n4477 2.71236
R8347 VSS.n4481 VSS.n4478 2.71236
R8348 VSS.n4489 VSS.n4454 2.71236
R8349 VSS.n4491 VSS.n4490 2.71236
R8350 VSS.n1999 VSS.n1998 2.71236
R8351 VSS.n2022 VSS.n2021 2.71236
R8352 VSS.n4359 VSS.n2023 2.71236
R8353 VSS.n4358 VSS.n4355 2.71236
R8354 VSS.n4354 VSS.n2024 2.71236
R8355 VSS.n4351 VSS.n4350 2.71236
R8356 VSS.n2031 VSS.n2025 2.71236
R8357 VSS.n4344 VSS.n2034 2.71236
R8358 VSS.n4343 VSS.n4341 2.71236
R8359 VSS.n4340 VSS.n4339 2.71236
R8360 VSS.n4113 VSS.n13 2.64083
R8361 VSS.n4788 VSS.n4787 2.64083
R8362 VSS.n4133 VSS.n4132 2.61497
R8363 VSS.n4192 VSS.n4073 2.61497
R8364 VSS.n493 VSS.n483 2.61497
R8365 VSS.n5230 VSS.n313 2.61497
R8366 VSS.n5276 VSS.n294 2.61497
R8367 VSS.n5322 VSS.n275 2.61497
R8368 VSS.n4789 VSS.n1215 2.61497
R8369 VSS.n4204 VSS.n4073 2.61359
R8370 VSS.n2693 VSS.n2659 2.60389
R8371 VSS.n3062 VSS.n2746 2.60389
R8372 VSS.n3027 VSS.n2809 2.60389
R8373 VSS.n4493 VSS.n4492 2.60389
R8374 VSS.n4320 VSS.n2053 2.60389
R8375 VSS.n4012 VSS.n4011 2.59839
R8376 VSS.n3189 VSS.n3188 2.59839
R8377 VSS.n3421 VSS.n3420 2.59839
R8378 VSS.n3000 VSS.n2927 2.59839
R8379 VSS.n4523 VSS.n1667 2.59839
R8380 VSS.n5414 VSS.n127 2.59839
R8381 VSS.n5121 VSS.n162 2.59839
R8382 VSS.n5053 VSS.n662 2.59839
R8383 VSS.n4893 VSS.n675 2.59839
R8384 VSS.n4738 VSS.n868 2.59839
R8385 VSS.n4140 VSS.n4089 2.58636
R8386 VSS.n1488 VSS.n1406 2.45707
R8387 VSS.n4222 VSS.n4221 2.45707
R8388 VSS.n4013 VSS.n2078 2.45707
R8389 VSS.n4683 VSS.n4650 2.45707
R8390 VSS.n4259 VSS.n4253 2.3255
R8391 VSS.n4261 VSS.n4260 2.3255
R8392 VSS.n497 VSS.n483 2.28816
R8393 VSS.n5231 VSS.n5230 2.28816
R8394 VSS.n5277 VSS.n5276 2.28816
R8395 VSS.n5323 VSS.n5322 2.28816
R8396 VSS.n4793 VSS.n1215 2.28816
R8397 VSS.n3101 VSS.n2659 2.27847
R8398 VSS.n3066 VSS.n2746 2.27847
R8399 VSS.n3031 VSS.n2809 2.27847
R8400 VSS.n4492 VSS.n4491 2.27847
R8401 VSS.n4339 VSS.n2053 2.27847
R8402 VSS.n3124 VSS.n2584 2.16999
R8403 VSS.n3123 VSS.n2585 2.16999
R8404 VSS.n2633 VSS.n2630 2.16999
R8405 VSS.n3117 VSS.n3116 2.16999
R8406 VSS.n3113 VSS.n2634 2.16999
R8407 VSS.n3112 VSS.n2635 2.16999
R8408 VSS.n2642 VSS.n2639 2.16999
R8409 VSS.n3106 VSS.n3105 2.16999
R8410 VSS.n3103 VSS.n3102 2.16999
R8411 VSS.n3092 VSS.n3091 2.16999
R8412 VSS.n3088 VSS.n2713 2.16999
R8413 VSS.n2720 VSS.n2717 2.16999
R8414 VSS.n3082 VSS.n3081 2.16999
R8415 VSS.n3078 VSS.n2721 2.16999
R8416 VSS.n3077 VSS.n2722 2.16999
R8417 VSS.n2729 VSS.n2726 2.16999
R8418 VSS.n3071 VSS.n3070 2.16999
R8419 VSS.n3068 VSS.n3067 2.16999
R8420 VSS.n2795 VSS.n2781 2.16999
R8421 VSS.n2797 VSS.n2796 2.16999
R8422 VSS.n3051 VSS.n3050 2.16999
R8423 VSS.n3047 VSS.n3046 2.16999
R8424 VSS.n3043 VSS.n2798 2.16999
R8425 VSS.n3042 VSS.n2799 2.16999
R8426 VSS.n2808 VSS.n2805 2.16999
R8427 VSS.n3036 VSS.n3035 2.16999
R8428 VSS.n3033 VSS.n3032 2.16999
R8429 VSS.n4633 VSS.n4632 2.16999
R8430 VSS.n4461 VSS.n1759 2.16999
R8431 VSS.n4462 VSS.n4460 2.16999
R8432 VSS.n4472 VSS.n4471 2.16999
R8433 VSS.n4475 VSS.n4458 2.16999
R8434 VSS.n4477 VSS.n4476 2.16999
R8435 VSS.n4482 VSS.n4481 2.16999
R8436 VSS.n4478 VSS.n4454 2.16999
R8437 VSS.n4490 VSS.n4489 2.16999
R8438 VSS.n2021 VSS.n2002 2.16999
R8439 VSS.n2023 VSS.n2022 2.16999
R8440 VSS.n4359 VSS.n4358 2.16999
R8441 VSS.n4355 VSS.n4354 2.16999
R8442 VSS.n4351 VSS.n2024 2.16999
R8443 VSS.n4350 VSS.n2025 2.16999
R8444 VSS.n2034 VSS.n2031 2.16999
R8445 VSS.n4344 VSS.n4343 2.16999
R8446 VSS.n4341 VSS.n4340 2.16999
R8447 VSS.n3965 VSS.n2170 2.12075
R8448 VSS.n3958 VSS.n2217 2.12075
R8449 VSS.n1891 VSS.n1889 2.12075
R8450 VSS.n3445 VSS.n2325 2.12075
R8451 VSS.n5497 VSS.n11 2.07029
R8452 VSS.n5193 VSS.n330 2.07029
R8453 VSS.n5239 VSS.n309 2.07029
R8454 VSS.n5285 VSS.n290 2.07029
R8455 VSS.n1204 VSS.n1203 2.07029
R8456 VSS.n2584 VSS.n2583 2.06152
R8457 VSS.n3093 VSS.n3092 2.06152
R8458 VSS.n2781 VSS.n2779 2.06152
R8459 VSS.n4634 VSS.n4633 2.06152
R8460 VSS.n2005 VSS.n2002 2.06152
R8461 VSS.n4271 VSS.n4239 1.89388
R8462 VSS.n4244 VSS.n4243 1.86266
R8463 VSS.n4245 VSS.n4240 1.8605
R8464 VSS.n4289 VSS.n4288 1.8605
R8465 VSS.n3965 VSS.n3964 1.8459
R8466 VSS.n3956 VSS.n2217 1.8459
R8467 VSS.n4562 VSS.n1891 1.8459
R8468 VSS.n3445 VSS.n3444 1.8459
R8469 VSS.n4781 VSS.n4780 1.80664
R8470 VSS.n1535 VSS.n1381 1.77399
R8471 VSS.n2114 VSS.n2068 1.76337
R8472 VSS.n1510 VSS.n1509 1.76337
R8473 VSS.n1556 VSS.n1537 1.61978
R8474 VSS.n4318 VSS.n4317 1.52394
R8475 VSS.n4286 VSS.n4285 1.52394
R8476 VSS.n4300 VSS.n4299 1.52302
R8477 VSS.n1509 VSS.n1322 1.45679
R8478 VSS.n4132 VSS.n18 1.41667
R8479 VSS.n4011 VSS.n4010 1.40769
R8480 VSS.n3193 VSS.n3189 1.40769
R8481 VSS.n3422 VSS.n3421 1.40769
R8482 VSS.n2927 VSS.n2926 1.40769
R8483 VSS.n4708 VSS.n1667 1.40769
R8484 VSS.n5415 VSS.n5414 1.40769
R8485 VSS.n5122 VSS.n5121 1.40769
R8486 VSS.n2423 VSS.n662 1.40769
R8487 VSS.n4894 VSS.n4893 1.40769
R8488 VSS.n4743 VSS.n4738 1.40769
R8489 VSS.n4192 VSS.n4191 1.38944
R8490 VSS.n3188 VSS.n2494 1.38063
R8491 VSS.n3420 VSS.n2459 1.38063
R8492 VSS.n3000 VSS.n2906 1.38063
R8493 VSS.n4523 VSS.n1989 1.38063
R8494 VSS.n162 VSS.n159 1.38063
R8495 VSS.n5053 VSS.n659 1.38063
R8496 VSS.n675 VSS.n673 1.38063
R8497 VSS.n868 VSS.n865 1.38063
R8498 VSS.n3154 VSS.n2494 1.35357
R8499 VSS.n3386 VSS.n2459 1.35357
R8500 VSS.n2906 VSS.n2903 1.35357
R8501 VSS.n1989 VSS.n1965 1.35357
R8502 VSS.n5379 VSS.n159 1.35357
R8503 VSS.n5086 VSS.n659 1.35357
R8504 VSS.n5049 VSS.n673 1.35357
R8505 VSS.n4858 VSS.n865 1.35357
R8506 VSS.n3152 VSS.n3151 1.29944
R8507 VSS.n3384 VSS.n3383 1.29944
R8508 VSS.n2902 VSS.n2901 1.29944
R8509 VSS.n4434 VSS.n4433 1.29944
R8510 VSS.n4685 VSS.n1726 1.29944
R8511 VSS.n5380 VSS.n151 1.29944
R8512 VSS.n5087 VSS.n651 1.29944
R8513 VSS.n3511 VSS.n670 1.29944
R8514 VSS.n4859 VSS.n858 1.29944
R8515 VSS.n1480 VSS.n1407 1.29944
R8516 VSS.n1010 VSS.n1009 1.29343
R8517 VSS.n3643 VSS.n3642 1.29343
R8518 VSS.n5001 VSS.n5000 1.29343
R8519 VSS.n267 VSS.n266 1.29343
R8520 VSS.n2202 VSS.n159 1.22878
R8521 VSS.n3930 VSS.n659 1.22878
R8522 VSS.n4556 VSS.n865 1.22878
R8523 VSS.n2941 VSS.n673 1.22878
R8524 VSS.n4518 VSS.n1989 1.22878
R8525 VSS.n2755 VSS.n2459 1.22878
R8526 VSS.n2906 VSS.n2817 1.22878
R8527 VSS.n2676 VSS.n2494 1.22878
R8528 VSS.n524 VSS.n523 1.14433
R8529 VSS.n567 VSS.n566 1.14433
R8530 VSS.n3802 VSS.n3630 1.14433
R8531 VSS.n1581 VSS.n1320 1.14433
R8532 VSS.n1560 VSS.n1341 1.14433
R8533 VSS.n1174 VSS.n1173 1.14433
R8534 VSS.n1153 VSS.n1152 1.14433
R8535 VSS.n3600 VSS.n2302 1.14433
R8536 VSS.n3567 VSS.n3566 1.14433
R8537 VSS.n3781 VSS.n3780 1.14433
R8538 VSS.n3313 VSS.n3308 1.13948
R8539 VSS.n3967 VSS.n3966 1.13948
R8540 VSS.n4566 VSS.n1886 1.13948
R8541 VSS.n3446 VSS.n2323 1.13948
R8542 VSS.n4778 VSS.n1254 1.13948
R8543 VSS.n3151 VSS.n3150 1.13708
R8544 VSS.n3383 VSS.n3382 1.13708
R8545 VSS.n2901 VSS.n2900 1.13708
R8546 VSS.n4434 VSS.n4432 1.13708
R8547 VSS.n1818 VSS.n1726 1.13708
R8548 VSS.n5384 VSS.n151 1.13708
R8549 VSS.n5091 VSS.n651 1.13708
R8550 VSS.n3511 VSS.n3510 1.13708
R8551 VSS.n4863 VSS.n858 1.13708
R8552 VSS.n1481 VSS.n1480 1.13708
R8553 VSS.n5476 VSS.n20 1.08986
R8554 VSS.n24 VSS.n21 1.08986
R8555 VSS.n5471 VSS.n25 1.08986
R8556 VSS.n33 VSS.n28 1.08986
R8557 VSS.n5465 VSS.n5464 1.08986
R8558 VSS.n462 VSS.n39 1.08986
R8559 VSS.n471 VSS.n470 1.08986
R8560 VSS.n518 VSS.n517 1.08986
R8561 VSS.n5455 VSS.n62 1.08986
R8562 VSS.n66 VSS.n63 1.08986
R8563 VSS.n5450 VSS.n67 1.08986
R8564 VSS.n75 VSS.n70 1.08986
R8565 VSS.n5444 VSS.n5443 1.08986
R8566 VSS.n553 VSS.n78 1.08986
R8567 VSS.n556 VSS.n551 1.08986
R8568 VSS.n561 VSS.n560 1.08986
R8569 VSS.n5175 VSS.n337 1.08986
R8570 VSS.n5171 VSS.n5170 1.08986
R8571 VSS.n5166 VSS.n342 1.08986
R8572 VSS.n3684 VSS.n343 1.08986
R8573 VSS.n3688 VSS.n3682 1.08986
R8574 VSS.n3707 VSS.n3675 1.08986
R8575 VSS.n3702 VSS.n3673 1.08986
R8576 VSS.n3730 VSS.n3672 1.08986
R8577 VSS.n4836 VSS.n4835 1.08986
R8578 VSS.n1298 VSS.n1295 1.08986
R8579 VSS.n1611 VSS.n1297 1.08986
R8580 VSS.n1601 VSS.n1301 1.08986
R8581 VSS.n1605 VSS.n1604 1.08986
R8582 VSS.n1596 VSS.n1310 1.08986
R8583 VSS.n1586 VSS.n1314 1.08986
R8584 VSS.n1590 VSS.n1589 1.08986
R8585 VSS.n1182 VSS.n912 1.08986
R8586 VSS.n4829 VSS.n913 1.08986
R8587 VSS.n4825 VSS.n4824 1.08986
R8588 VSS.n1356 VSS.n1355 1.08986
R8589 VSS.n1360 VSS.n1352 1.08986
R8590 VSS.n1369 VSS.n1346 1.08986
R8591 VSS.n1373 VSS.n1345 1.08986
R8592 VSS.n1378 VSS.n1342 1.08986
R8593 VSS.n4957 VSS.n720 1.08986
R8594 VSS.n4962 VSS.n4961 1.08986
R8595 VSS.n1049 VSS.n1048 1.08986
R8596 VSS.n1055 VSS.n1054 1.08986
R8597 VSS.n1068 VSS.n1045 1.08986
R8598 VSS.n1074 VSS.n1041 1.08986
R8599 VSS.n1079 VSS.n1078 1.08986
R8600 VSS.n1084 VSS.n1083 1.08986
R8601 VSS.n4932 VSS.n747 1.08986
R8602 VSS.n751 VSS.n748 1.08986
R8603 VSS.n4927 VSS.n753 1.08986
R8604 VSS.n4923 VSS.n4922 1.08986
R8605 VSS.n4919 VSS.n761 1.08986
R8606 VSS.n1138 VSS.n1137 1.08986
R8607 VSS.n1143 VSS.n1142 1.08986
R8608 VSS.n1147 VSS.n1146 1.08986
R8609 VSS.n3810 VSS.n2275 1.08986
R8610 VSS.n3844 VSS.n2276 1.08986
R8611 VSS.n3833 VSS.n2279 1.08986
R8612 VSS.n3838 VSS.n3837 1.08986
R8613 VSS.n3628 VSS.n2284 1.08986
R8614 VSS.n3619 VSS.n2287 1.08986
R8615 VSS.n3615 VSS.n3614 1.08986
R8616 VSS.n3608 VSS.n2297 1.08986
R8617 VSS.n2267 VSS.n2257 1.08986
R8618 VSS.n3879 VSS.n2258 1.08986
R8619 VSS.n3868 VSS.n2261 1.08986
R8620 VSS.n3873 VSS.n3872 1.08986
R8621 VSS.n3539 VSS.n3538 1.08986
R8622 VSS.n3554 VSS.n2315 1.08986
R8623 VSS.n2316 VSS.n2312 1.08986
R8624 VSS.n3561 VSS.n3560 1.08986
R8625 VSS.n5160 VSS.n365 1.08986
R8626 VSS.n369 VSS.n366 1.08986
R8627 VSS.n5155 VSS.n371 1.08986
R8628 VSS.n5151 VSS.n5150 1.08986
R8629 VSS.n5147 VSS.n376 1.08986
R8630 VSS.n3766 VSS.n3765 1.08986
R8631 VSS.n3771 VSS.n3770 1.08986
R8632 VSS.n3775 VSS.n3774 1.08986
R8633 VSS.n3204 VSS.n3201 1.08525
R8634 VSS.n3343 VSS.n3202 1.08525
R8635 VSS.n3212 VSS.n3208 1.08525
R8636 VSS.n3337 VSS.n3336 1.08525
R8637 VSS.n3333 VSS.n3215 1.08525
R8638 VSS.n3324 VSS.n3220 1.08525
R8639 VSS.n3320 VSS.n3319 1.08525
R8640 VSS.n3231 VSS.n3228 1.08525
R8641 VSS.n3997 VSS.n2117 1.08525
R8642 VSS.n3993 VSS.n3992 1.08525
R8643 VSS.n3989 VSS.n2124 1.08525
R8644 VSS.n2126 VSS.n2125 1.08525
R8645 VSS.n3984 VSS.n2129 1.08525
R8646 VSS.n3976 VSS.n2139 1.08525
R8647 VSS.n3973 VSS.n2141 1.08525
R8648 VSS.n2147 VSS.n2145 1.08525
R8649 VSS.n2326 VSS.n1838 1.08525
R8650 VSS.n4596 VSS.n1839 1.08525
R8651 VSS.n1848 VSS.n1843 1.08525
R8652 VSS.n4590 VSS.n4589 1.08525
R8653 VSS.n4586 VSS.n1851 1.08525
R8654 VSS.n4577 VSS.n1856 1.08525
R8655 VSS.n4573 VSS.n4572 1.08525
R8656 VSS.n1867 VSS.n1864 1.08525
R8657 VSS.n2223 VSS.n2218 1.08525
R8658 VSS.n3916 VSS.n3915 1.08525
R8659 VSS.n2353 VSS.n2352 1.08525
R8660 VSS.n2358 VSS.n2357 1.08525
R8661 VSS.n2362 VSS.n2361 1.08525
R8662 VSS.n2371 VSS.n2341 1.08525
R8663 VSS.n2375 VSS.n2343 1.08525
R8664 VSS.n3438 VSS.n3437 1.08525
R8665 VSS.n4719 VSS.n1621 1.08525
R8666 VSS.n1895 VSS.n1622 1.08525
R8667 VSS.n1898 VSS.n1892 1.08525
R8668 VSS.n1941 VSS.n1940 1.08525
R8669 VSS.n1937 VSS.n1902 1.08525
R8670 VSS.n1907 VSS.n1905 1.08525
R8671 VSS.n1927 VSS.n1926 1.08525
R8672 VSS.n1920 VSS.n1919 1.08525
R8673 VSS.n4009 VSS.n4006 1.08295
R8674 VSS.n2535 VSS.n2534 1.08295
R8675 VSS.n2540 VSS.n2539 1.08295
R8676 VSS.n2574 VSS.n2543 1.08295
R8677 VSS.n2570 VSS.n2569 1.08295
R8678 VSS.n2552 VSS.n2551 1.08295
R8679 VSS.n2561 VSS.n2555 1.08295
R8680 VSS.n2557 VSS.n2518 1.08295
R8681 VSS.n3192 VSS.n2487 1.08295
R8682 VSS.n3373 VSS.n2488 1.08295
R8683 VSS.n3369 VSS.n3368 1.08295
R8684 VSS.n3244 VSS.n3243 1.08295
R8685 VSS.n3248 VSS.n3242 1.08295
R8686 VSS.n3257 VSS.n3236 1.08295
R8687 VSS.n3268 VSS.n3262 1.08295
R8688 VSS.n3266 VSS.n2466 1.08295
R8689 VSS.n3432 VSS.n2395 1.08295
R8690 VSS.n2399 VSS.n2396 1.08295
R8691 VSS.n2869 VSS.n2866 1.08295
R8692 VSS.n2871 VSS.n2862 1.08295
R8693 VSS.n2875 VSS.n2861 1.08295
R8694 VSS.n2884 VSS.n2857 1.08295
R8695 VSS.n2889 VSS.n2854 1.08295
R8696 VSS.n2893 VSS.n2853 1.08295
R8697 VSS.n2925 VSS.n1780 1.08295
R8698 VSS.n4626 VSS.n1781 1.08295
R8699 VSS.n4622 VSS.n4621 1.08295
R8700 VSS.n4403 VSS.n4402 1.08295
R8701 VSS.n4407 VSS.n4401 1.08295
R8702 VSS.n4416 VSS.n4370 1.08295
R8703 VSS.n4421 VSS.n4369 1.08295
R8704 VSS.n4425 VSS.n4368 1.08295
R8705 VSS.n4690 VSS.n1669 1.08295
R8706 VSS.n4714 VSS.n1644 1.08295
R8707 VSS.n1789 VSS.n1645 1.08295
R8708 VSS.n1795 VSS.n1792 1.08295
R8709 VSS.n1797 VSS.n1788 1.08295
R8710 VSS.n1808 VSS.n1787 1.08295
R8711 VSS.n1815 VSS.n1813 1.08295
R8712 VSS.n1823 VSS.n1822 1.08295
R8713 VSS.n5435 VSS.n101 1.08295
R8714 VSS.n105 VSS.n102 1.08295
R8715 VSS.n5406 VSS.n5405 1.08295
R8716 VSS.n5402 VSS.n133 1.08295
R8717 VSS.n135 VSS.n134 1.08295
R8718 VSS.n5393 VSS.n5392 1.08295
R8719 VSS.n5389 VSS.n148 1.08295
R8720 VSS.n150 VSS.n149 1.08295
R8721 VSS.n5142 VSS.n397 1.08295
R8722 VSS.n401 VSS.n398 1.08295
R8723 VSS.n5113 VSS.n5112 1.08295
R8724 VSS.n5109 VSS.n633 1.08295
R8725 VSS.n635 VSS.n634 1.08295
R8726 VSS.n5100 VSS.n5099 1.08295
R8727 VSS.n5096 VSS.n648 1.08295
R8728 VSS.n650 VSS.n649 1.08295
R8729 VSS.n2422 VSS.n2243 1.08295
R8730 VSS.n3909 VSS.n2244 1.08295
R8731 VSS.n3905 VSS.n3904 1.08295
R8732 VSS.n3474 VSS.n3473 1.08295
R8733 VSS.n3478 VSS.n3472 1.08295
R8734 VSS.n3489 VSS.n3468 1.08295
R8735 VSS.n3500 VSS.n3467 1.08295
R8736 VSS.n3505 VSS.n3504 1.08295
R8737 VSS.n4914 VSS.n782 1.08295
R8738 VSS.n786 VSS.n783 1.08295
R8739 VSS.n4885 VSS.n4884 1.08295
R8740 VSS.n4881 VSS.n840 1.08295
R8741 VSS.n842 VSS.n841 1.08295
R8742 VSS.n4872 VSS.n4871 1.08295
R8743 VSS.n4868 VSS.n855 1.08295
R8744 VSS.n857 VSS.n856 1.08295
R8745 VSS.n4742 VSS.n1276 1.08295
R8746 VSS.n4771 VSS.n1277 1.08295
R8747 VSS.n4767 VSS.n4766 1.08295
R8748 VSS.n1418 VSS.n1417 1.08295
R8749 VSS.n1422 VSS.n1414 1.08295
R8750 VSS.n1440 VSS.n1412 1.08295
R8751 VSS.n1445 VSS.n1411 1.08295
R8752 VSS.n1448 VSS.n1410 1.08295
R8753 VSS.n5460 VSS 1.06263
R8754 VSS.n5440 VSS 1.06263
R8755 VSS VSS.n3693 1.06263
R8756 VSS VSS.n1307 1.06263
R8757 VSS VSS.n1350 1.06263
R8758 VSS VSS.n1042 1.06263
R8759 VSS.n1134 VSS 1.06263
R8760 VSS VSS.n2286 1.06263
R8761 VSS.n3548 VSS 1.06263
R8762 VSS.n3762 VSS 1.06263
R8763 VSS VSS.n3217 1.05813
R8764 VSS VSS.n3979 1.05813
R8765 VSS VSS.n1853 1.05813
R8766 VSS.n2369 VSS 1.05813
R8767 VSS.n1910 VSS 1.05813
R8768 VSS.n2566 VSS 1.05589
R8769 VSS VSS.n3237 1.05589
R8770 VSS VSS.n2858 1.05589
R8771 VSS VSS.n4371 1.05589
R8772 VSS.n1806 VSS 1.05589
R8773 VSS.n143 VSS 1.05589
R8774 VSS.n643 VSS 1.05589
R8775 VSS.n3494 VSS 1.05589
R8776 VSS.n850 VSS 1.05589
R8777 VSS.n1437 VSS 1.05589
R8778 VSS.n20 VSS.n18 1.03539
R8779 VSS.n4190 VSS.n62 1.03539
R8780 VSS.n5176 VSS.n5175 1.03539
R8781 VSS.n4836 VSS.n890 1.03539
R8782 VSS.n1183 VSS.n1182 1.03539
R8783 VSS.n4938 VSS.n720 1.03539
R8784 VSS.n820 VSS.n747 1.03539
R8785 VSS.n3811 VSS.n3810 1.03539
R8786 VSS.n2268 VSS.n2267 1.03539
R8787 VSS.n612 VSS.n365 1.03539
R8788 VSS.n3204 VSS.n2169 1.03101
R8789 VSS.n3998 VSS.n3997 1.03101
R8790 VSS.n2326 VSS.n2324 1.03101
R8791 VSS.n2441 VSS.n2218 1.03101
R8792 VSS.n1621 VSS.n1620 1.03101
R8793 VSS.n4010 VSS.n4009 1.02883
R8794 VSS.n3193 VSS.n3192 1.02883
R8795 VSS.n3422 VSS.n2395 1.02883
R8796 VSS.n2926 VSS.n2925 1.02883
R8797 VSS.n4708 VSS.n4690 1.02883
R8798 VSS.n5415 VSS.n101 1.02883
R8799 VSS.n5122 VSS.n397 1.02883
R8800 VSS.n2423 VSS.n2422 1.02883
R8801 VSS.n4894 VSS.n782 1.02883
R8802 VSS.n4743 VSS.n4742 1.02883
R8803 VSS.n4234 VSS.n4233 1.00976
R8804 VSS.n4235 VSS.n4234 1.00976
R8805 VSS.n524 VSS.n231 0.980926
R8806 VSS.n611 VSS.n567 0.980926
R8807 VSS.n5176 VSS.n231 0.980926
R8808 VSS.n3807 VSS.n3630 0.980926
R8809 VSS.n890 VSS.n887 0.980926
R8810 VSS.n1581 VSS.n1322 0.980926
R8811 VSS.n1183 VSS.n954 0.980926
R8812 VSS.n1537 VSS.n1341 0.980926
R8813 VSS.n4938 VSS.n719 0.980926
R8814 VSS.n1173 VSS.n954 0.980926
R8815 VSS.n820 VSS.n694 0.980926
R8816 VSS.n1153 VSS.n887 0.980926
R8817 VSS.n3811 VSS.n3807 0.980926
R8818 VSS.n3600 VSS.n719 0.980926
R8819 VSS.n2268 VSS.n192 0.980926
R8820 VSS.n3567 VSS.n694 0.980926
R8821 VSS.n612 VSS.n611 0.980926
R8822 VSS.n3781 VSS.n192 0.980926
R8823 VSS.n3965 VSS.n2169 0.976771
R8824 VSS.n3308 VSS.n2217 0.976771
R8825 VSS.n3998 VSS.n2115 0.976771
R8826 VSS.n3966 VSS.n3965 0.976771
R8827 VSS.n3445 VSS.n2324 0.976771
R8828 VSS.n1891 VSS.n1886 0.976771
R8829 VSS.n2441 VSS.n2217 0.976771
R8830 VSS.n3446 VSS.n3445 0.976771
R8831 VSS.n1891 VSS.n1620 0.976771
R8832 VSS.n4779 VSS.n4778 0.976771
R8833 VSS.n5476 VSS.n5475 0.926457
R8834 VSS.n5472 VSS.n24 0.926457
R8835 VSS.n44 VSS.n25 0.926457
R8836 VSS.n33 VSS.n31 0.926457
R8837 VSS.n5464 VSS.n32 0.926457
R8838 VSS.n5460 VSS.n5459 0.926457
R8839 VSS.n463 VSS.n462 0.926457
R8840 VSS.n471 VSS.n461 0.926457
R8841 VSS.n517 VSS.n459 0.926457
R8842 VSS.n5455 VSS.n5454 0.926457
R8843 VSS.n5451 VSS.n66 0.926457
R8844 VSS.n83 VSS.n67 0.926457
R8845 VSS.n76 VSS.n75 0.926457
R8846 VSS.n5443 VSS.n77 0.926457
R8847 VSS.n5440 VSS.n5439 0.926457
R8848 VSS.n553 VSS.n552 0.926457
R8849 VSS.n557 VSS.n556 0.926457
R8850 VSS.n560 VSS.n543 0.926457
R8851 VSS.n339 VSS.n337 0.926457
R8852 VSS.n5170 VSS.n340 0.926457
R8853 VSS.n5166 VSS.n5165 0.926457
R8854 VSS.n3684 VSS.n3683 0.926457
R8855 VSS.n3689 VSS.n3688 0.926457
R8856 VSS.n3693 VSS.n3692 0.926457
R8857 VSS.n3707 VSS.n3706 0.926457
R8858 VSS.n3703 VSS.n3673 0.926457
R8859 VSS.n3801 VSS.n3730 0.926457
R8860 VSS.n4835 VSS.n891 0.926457
R8861 VSS.n1612 VSS.n1295 0.926457
R8862 VSS.n1303 VSS.n1297 0.926457
R8863 VSS.n1601 VSS.n1306 0.926457
R8864 VSS.n1604 VSS.n1600 0.926457
R8865 VSS.n1597 VSS.n1307 0.926457
R8866 VSS.n1316 VSS.n1310 0.926457
R8867 VSS.n1586 VSS.n1319 0.926457
R8868 VSS.n1589 VSS.n1585 0.926457
R8869 VSS.n4830 VSS.n912 0.926457
R8870 VSS.n916 VSS.n913 0.926457
R8871 VSS.n4824 VSS.n917 0.926457
R8872 VSS.n1359 VSS.n1356 0.926457
R8873 VSS.n1365 VSS.n1352 0.926457
R8874 VSS.n1368 VSS.n1350 0.926457
R8875 VSS.n1374 VSS.n1346 0.926457
R8876 VSS.n1377 VSS.n1345 0.926457
R8877 VSS.n1561 VSS.n1342 0.926457
R8878 VSS.n4957 VSS.n722 0.926457
R8879 VSS.n4961 VSS.n723 0.926457
R8880 VSS.n1050 VSS.n1049 0.926457
R8881 VSS.n1054 VSS.n1053 0.926457
R8882 VSS.n1068 VSS.n1067 0.926457
R8883 VSS.n1064 VSS.n1042 0.926457
R8884 VSS.n1077 VSS.n1074 0.926457
R8885 VSS.n1078 VSS.n1039 0.926457
R8886 VSS.n1084 VSS.n1036 0.926457
R8887 VSS.n4932 VSS.n4931 0.926457
R8888 VSS.n4928 VSS.n751 0.926457
R8889 VSS.n759 VSS.n753 0.926457
R8890 VSS.n4922 VSS.n760 0.926457
R8891 VSS.n4919 VSS.n4918 0.926457
R8892 VSS.n1134 VSS.n1129 0.926457
R8893 VSS.n1137 VSS.n1127 0.926457
R8894 VSS.n1143 VSS.n1125 0.926457
R8895 VSS.n1146 VSS.n1123 0.926457
R8896 VSS.n3845 VSS.n2275 0.926457
R8897 VSS.n2278 VSS.n2276 0.926457
R8898 VSS.n3833 VSS.n2281 0.926457
R8899 VSS.n3837 VSS.n2282 0.926457
R8900 VSS.n3628 VSS.n3627 0.926457
R8901 VSS.n3620 VSS.n2286 0.926457
R8902 VSS.n2294 VSS.n2287 0.926457
R8903 VSS.n3614 VSS.n2295 0.926457
R8904 VSS.n3608 VSS.n3607 0.926457
R8905 VSS.n3880 VSS.n2257 0.926457
R8906 VSS.n2260 VSS.n2258 0.926457
R8907 VSS.n3868 VSS.n2263 0.926457
R8908 VSS.n3872 VSS.n2264 0.926457
R8909 VSS.n3538 VSS.n3537 0.926457
R8910 VSS.n3549 VSS.n3548 0.926457
R8911 VSS.n3554 VSS.n3553 0.926457
R8912 VSS.n2312 VSS.n2311 0.926457
R8913 VSS.n3560 VSS.n2309 0.926457
R8914 VSS.n5160 VSS.n5159 0.926457
R8915 VSS.n5156 VSS.n369 0.926457
R8916 VSS.n374 VSS.n371 0.926457
R8917 VSS.n5150 VSS.n375 0.926457
R8918 VSS.n5147 VSS.n5146 0.926457
R8919 VSS.n3762 VSS.n3757 0.926457
R8920 VSS.n3765 VSS.n3755 0.926457
R8921 VSS.n3771 VSS.n3753 0.926457
R8922 VSS.n3774 VSS.n3751 0.926457
R8923 VSS.n3344 VSS.n3201 0.922534
R8924 VSS.n3207 VSS.n3202 0.922534
R8925 VSS.n3213 VSS.n3212 0.922534
R8926 VSS.n3336 VSS.n3214 0.922534
R8927 VSS.n3333 VSS.n3332 0.922534
R8928 VSS.n3325 VSS.n3217 0.922534
R8929 VSS.n3227 VSS.n3220 0.922534
R8930 VSS.n3319 VSS.n3317 0.922534
R8931 VSS.n3314 VSS.n3231 0.922534
R8932 VSS.n2120 VSS.n2117 0.922534
R8933 VSS.n3992 VSS.n2123 0.922534
R8934 VSS.n3989 VSS.n3988 0.922534
R8935 VSS.n3985 VSS.n2126 0.922534
R8936 VSS.n2135 VSS.n2129 0.922534
R8937 VSS.n3979 VSS.n2138 0.922534
R8938 VSS.n3976 VSS.n3975 0.922534
R8939 VSS.n2144 VSS.n2141 0.922534
R8940 VSS.n2149 VSS.n2147 0.922534
R8941 VSS.n4597 VSS.n1838 0.922534
R8942 VSS.n1842 VSS.n1839 0.922534
R8943 VSS.n1849 VSS.n1848 0.922534
R8944 VSS.n4589 VSS.n1850 0.922534
R8945 VSS.n4586 VSS.n4585 0.922534
R8946 VSS.n4578 VSS.n1853 0.922534
R8947 VSS.n1863 VSS.n1856 0.922534
R8948 VSS.n4572 VSS.n4570 0.922534
R8949 VSS.n4567 VSS.n1867 0.922534
R8950 VSS.n2223 VSS.n2220 0.922534
R8951 VSS.n3915 VSS.n2221 0.922534
R8952 VSS.n2352 VSS.n2351 0.922534
R8953 VSS.n2358 VSS.n2346 0.922534
R8954 VSS.n2361 VSS.n2348 0.922534
R8955 VSS.n2370 VSS.n2369 0.922534
R8956 VSS.n2376 VSS.n2341 0.922534
R8957 VSS.n2343 VSS.n2332 0.922534
R8958 VSS.n3437 VSS.n3436 0.922534
R8959 VSS.n4719 VSS.n4718 0.922534
R8960 VSS.n1895 VSS.n1894 0.922534
R8961 VSS.n1900 VSS.n1898 0.922534
R8962 VSS.n1940 VSS.n1901 0.922534
R8963 VSS.n1937 VSS.n1936 0.922534
R8964 VSS.n1911 VSS.n1910 0.922534
R8965 VSS.n1914 VSS.n1907 0.922534
R8966 VSS.n1926 VSS.n1924 0.922534
R8967 VSS.n1921 VSS.n1920 0.922534
R8968 VSS.n4006 VSS.n2083 0.920585
R8969 VSS.n2534 VSS.n2533 0.920585
R8970 VSS.n2575 VSS.n2540 0.920585
R8971 VSS.n2544 VSS.n2543 0.920585
R8972 VSS.n2569 VSS.n2546 0.920585
R8973 VSS.n2566 VSS.n2565 0.920585
R8974 VSS.n2562 VSS.n2552 0.920585
R8975 VSS.n2556 VSS.n2555 0.920585
R8976 VSS.n3147 VSS.n2518 0.920585
R8977 VSS.n3374 VSS.n2487 0.920585
R8978 VSS.n2489 VSS.n2488 0.920585
R8979 VSS.n3368 VSS.n2491 0.920585
R8980 VSS.n3249 VSS.n3243 0.920585
R8981 VSS.n3252 VSS.n3242 0.920585
R8982 VSS.n3258 VSS.n3237 0.920585
R8983 VSS.n3261 VSS.n3236 0.920585
R8984 VSS.n3268 VSS.n3267 0.920585
R8985 VSS.n3379 VSS.n2466 0.920585
R8986 VSS.n3432 VSS.n3431 0.920585
R8987 VSS.n2400 VSS.n2399 0.920585
R8988 VSS.n2870 VSS.n2869 0.920585
R8989 VSS.n2876 VSS.n2862 0.920585
R8990 VSS.n2879 VSS.n2861 0.920585
R8991 VSS.n2885 VSS.n2858 0.920585
R8992 VSS.n2888 VSS.n2857 0.920585
R8993 VSS.n2894 VSS.n2854 0.920585
R8994 VSS.n2897 VSS.n2853 0.920585
R8995 VSS.n4627 VSS.n1780 0.920585
R8996 VSS.n1827 VSS.n1781 0.920585
R8997 VSS.n4621 VSS.n1829 0.920585
R8998 VSS.n4408 VSS.n4402 0.920585
R8999 VSS.n4411 VSS.n4401 0.920585
R9000 VSS.n4417 VSS.n4371 0.920585
R9001 VSS.n4420 VSS.n4370 0.920585
R9002 VSS.n4426 VSS.n4369 0.920585
R9003 VSS.n4429 VSS.n4368 0.920585
R9004 VSS.n1669 VSS.n1668 0.920585
R9005 VSS.n4714 VSS.n4713 0.920585
R9006 VSS.n1790 VSS.n1789 0.920585
R9007 VSS.n1798 VSS.n1795 0.920585
R9008 VSS.n1801 VSS.n1788 0.920585
R9009 VSS.n1809 VSS.n1806 0.920585
R9010 VSS.n1812 VSS.n1787 0.920585
R9011 VSS.n1816 VSS.n1815 0.920585
R9012 VSS.n1822 VSS.n1821 0.920585
R9013 VSS.n5435 VSS.n5434 0.920585
R9014 VSS.n106 VSS.n105 0.920585
R9015 VSS.n5405 VSS.n132 0.920585
R9016 VSS.n5402 VSS.n5401 0.920585
R9017 VSS.n5398 VSS.n135 0.920585
R9018 VSS.n144 VSS.n143 0.920585
R9019 VSS.n5392 VSS.n147 0.920585
R9020 VSS.n5389 VSS.n5388 0.920585
R9021 VSS.n5385 VSS.n150 0.920585
R9022 VSS.n5142 VSS.n5141 0.920585
R9023 VSS.n402 VSS.n401 0.920585
R9024 VSS.n5112 VSS.n632 0.920585
R9025 VSS.n5109 VSS.n5108 0.920585
R9026 VSS.n5105 VSS.n635 0.920585
R9027 VSS.n644 VSS.n643 0.920585
R9028 VSS.n5099 VSS.n647 0.920585
R9029 VSS.n5096 VSS.n5095 0.920585
R9030 VSS.n5092 VSS.n650 0.920585
R9031 VSS.n3910 VSS.n2243 0.920585
R9032 VSS.n2247 VSS.n2244 0.920585
R9033 VSS.n3904 VSS.n2249 0.920585
R9034 VSS.n3479 VSS.n3473 0.920585
R9035 VSS.n3482 VSS.n3472 0.920585
R9036 VSS.n3494 VSS.n3493 0.920585
R9037 VSS.n3490 VSS.n3468 0.920585
R9038 VSS.n3503 VSS.n3500 0.920585
R9039 VSS.n3504 VSS.n3465 0.920585
R9040 VSS.n4914 VSS.n4913 0.920585
R9041 VSS.n787 VSS.n786 0.920585
R9042 VSS.n4884 VSS.n839 0.920585
R9043 VSS.n4881 VSS.n4880 0.920585
R9044 VSS.n4877 VSS.n842 0.920585
R9045 VSS.n851 VSS.n850 0.920585
R9046 VSS.n4871 VSS.n854 0.920585
R9047 VSS.n4868 VSS.n4867 0.920585
R9048 VSS.n4864 VSS.n857 0.920585
R9049 VSS.n4772 VSS.n1276 0.920585
R9050 VSS.n1280 VSS.n1277 0.920585
R9051 VSS.n4766 VSS.n1281 0.920585
R9052 VSS.n1421 VSS.n1418 0.920585
R9053 VSS.n1433 VSS.n1414 0.920585
R9054 VSS.n1437 VSS.n1436 0.920585
R9055 VSS.n1441 VSS.n1440 0.920585
R9056 VSS.n1445 VSS.n1444 0.920585
R9057 VSS.n1449 VSS.n1448 0.920585
R9058 VSS.n4841 VSS.n4840 0.903568
R9059 VSS.n958 VSS.n955 0.903568
R9060 VSS.n5032 VSS.n5031 0.903568
R9061 VSS.n5358 VSS.n5357 0.903568
R9062 VSS.n3631 VSS.n219 0.903568
R9063 VSS.n5011 VSS.n5010 0.903568
R9064 VSS.n5339 VSS.n5338 0.903568
R9065 VSS.n5362 VSS.n181 0.903568
R9066 VSS.n2208 VSS.n2170 0.903568
R9067 VSS.n3959 VSS.n3958 0.903568
R9068 VSS.n1954 VSS.n1889 0.903568
R9069 VSS.n2983 VSS.n2325 0.903568
R9070 VSS.n5504 VSS.n10 0.871989
R9071 VSS.n5505 VSS.n8 0.871989
R9072 VSS.n5510 VSS.n5509 0.871989
R9073 VSS.n5514 VSS.n4 0.871989
R9074 VSS.n5519 VSS.n1 0.871989
R9075 VSS.n488 VSS.n486 0.871989
R9076 VSS.n487 VSS.n482 0.871989
R9077 VSS.n498 VSS.n497 0.871989
R9078 VSS.n5200 VSS.n5198 0.871989
R9079 VSS.n5199 VSS.n326 0.871989
R9080 VSS.n5207 VSS.n5206 0.871989
R9081 VSS.n324 VSS.n323 0.871989
R9082 VSS.n5214 VSS.n321 0.871989
R9083 VSS.n5222 VSS.n5221 0.871989
R9084 VSS.n319 VSS.n318 0.871989
R9085 VSS.n5231 VSS.n315 0.871989
R9086 VSS.n5246 VSS.n5244 0.871989
R9087 VSS.n5245 VSS.n307 0.871989
R9088 VSS.n5253 VSS.n5252 0.871989
R9089 VSS.n305 VSS.n304 0.871989
R9090 VSS.n5260 VSS.n302 0.871989
R9091 VSS.n5268 VSS.n5267 0.871989
R9092 VSS.n300 VSS.n299 0.871989
R9093 VSS.n5277 VSS.n296 0.871989
R9094 VSS.n5292 VSS.n5290 0.871989
R9095 VSS.n5291 VSS.n288 0.871989
R9096 VSS.n5299 VSS.n5298 0.871989
R9097 VSS.n286 VSS.n285 0.871989
R9098 VSS.n5306 VSS.n283 0.871989
R9099 VSS.n5314 VSS.n5313 0.871989
R9100 VSS.n281 VSS.n280 0.871989
R9101 VSS.n5323 VSS.n277 0.871989
R9102 VSS.n4819 VSS.n4818 0.871989
R9103 VSS.n4814 VSS.n1205 0.871989
R9104 VSS.n4813 VSS.n4811 0.871989
R9105 VSS.n4810 VSS.n1209 0.871989
R9106 VSS.n4802 VSS.n1213 0.871989
R9107 VSS.n4801 VSS.n4798 0.871989
R9108 VSS.n4797 VSS.n1214 0.871989
R9109 VSS.n4794 VSS.n4793 0.871989
R9110 VSS.n1178 VSS.n954 0.82504
R9111 VSS.n3807 VSS.n3806 0.82504
R9112 VSS.n5008 VSS.n719 0.82504
R9113 VSS.n5336 VSS.n231 0.82504
R9114 VSS.n4840 VSS.n887 0.746512
R9115 VSS.n5031 VSS.n694 0.746512
R9116 VSS.n5357 VSS.n192 0.746512
R9117 VSS.n611 VSS.n181 0.746512
R9118 VSS.n4260 VSS.n4259 0.708416
R9119 VSS.n4306 VSS.n4236 0.699855
R9120 VSS.n4316 VSS 0.669484
R9121 VSS.n5515 VSS 0.599649
R9122 VSS VSS.n5213 0.599649
R9123 VSS VSS.n5259 0.599649
R9124 VSS VSS.n5305 0.599649
R9125 VSS.n4807 VSS 0.599649
R9126 VSS VSS.n4306 0.588917
R9127 VSS.n4301 VSS.n4300 0.52613
R9128 VSS.n4245 VSS.n4244 0.512067
R9129 VSS.n4299 VSS.n4298 0.506084
R9130 VSS VSS.n4246 0.450368
R9131 VSS.n5475 VSS.n21 0.436245
R9132 VSS.n5472 VSS.n5471 0.436245
R9133 VSS.n44 VSS.n28 0.436245
R9134 VSS.n5465 VSS.n31 0.436245
R9135 VSS.n5459 VSS.n39 0.436245
R9136 VSS.n470 VSS.n463 0.436245
R9137 VSS.n518 VSS.n461 0.436245
R9138 VSS.n523 VSS.n459 0.436245
R9139 VSS.n5454 VSS.n63 0.436245
R9140 VSS.n5451 VSS.n5450 0.436245
R9141 VSS.n83 VSS.n70 0.436245
R9142 VSS.n5444 VSS.n76 0.436245
R9143 VSS.n5439 VSS.n78 0.436245
R9144 VSS.n552 VSS.n551 0.436245
R9145 VSS.n561 VSS.n557 0.436245
R9146 VSS.n566 VSS.n543 0.436245
R9147 VSS.n5171 VSS.n339 0.436245
R9148 VSS.n342 VSS.n340 0.436245
R9149 VSS.n5165 VSS.n343 0.436245
R9150 VSS.n3683 VSS.n3682 0.436245
R9151 VSS.n3692 VSS.n3675 0.436245
R9152 VSS.n3706 VSS.n3702 0.436245
R9153 VSS.n3703 VSS.n3672 0.436245
R9154 VSS.n3802 VSS.n3801 0.436245
R9155 VSS.n1298 VSS.n891 0.436245
R9156 VSS.n1612 VSS.n1611 0.436245
R9157 VSS.n1303 VSS.n1301 0.436245
R9158 VSS.n1605 VSS.n1306 0.436245
R9159 VSS.n1597 VSS.n1596 0.436245
R9160 VSS.n1316 VSS.n1314 0.436245
R9161 VSS.n1590 VSS.n1319 0.436245
R9162 VSS.n1585 VSS.n1320 0.436245
R9163 VSS.n4830 VSS.n4829 0.436245
R9164 VSS.n4825 VSS.n916 0.436245
R9165 VSS.n1355 VSS.n917 0.436245
R9166 VSS.n1360 VSS.n1359 0.436245
R9167 VSS.n1369 VSS.n1368 0.436245
R9168 VSS.n1374 VSS.n1373 0.436245
R9169 VSS.n1378 VSS.n1377 0.436245
R9170 VSS.n1561 VSS.n1560 0.436245
R9171 VSS.n4962 VSS.n722 0.436245
R9172 VSS.n1048 VSS.n723 0.436245
R9173 VSS.n1055 VSS.n1050 0.436245
R9174 VSS.n1053 VSS.n1045 0.436245
R9175 VSS.n1064 VSS.n1041 0.436245
R9176 VSS.n1079 VSS.n1077 0.436245
R9177 VSS.n1083 VSS.n1039 0.436245
R9178 VSS.n1174 VSS.n1036 0.436245
R9179 VSS.n4931 VSS.n748 0.436245
R9180 VSS.n4928 VSS.n4927 0.436245
R9181 VSS.n4923 VSS.n759 0.436245
R9182 VSS.n761 VSS.n760 0.436245
R9183 VSS.n1138 VSS.n1129 0.436245
R9184 VSS.n1142 VSS.n1127 0.436245
R9185 VSS.n1147 VSS.n1125 0.436245
R9186 VSS.n1152 VSS.n1123 0.436245
R9187 VSS.n3845 VSS.n3844 0.436245
R9188 VSS.n2279 VSS.n2278 0.436245
R9189 VSS.n3838 VSS.n2281 0.436245
R9190 VSS.n2284 VSS.n2282 0.436245
R9191 VSS.n3620 VSS.n3619 0.436245
R9192 VSS.n3615 VSS.n2294 0.436245
R9193 VSS.n2297 VSS.n2295 0.436245
R9194 VSS.n3607 VSS.n2302 0.436245
R9195 VSS.n3880 VSS.n3879 0.436245
R9196 VSS.n2261 VSS.n2260 0.436245
R9197 VSS.n3873 VSS.n2263 0.436245
R9198 VSS.n3539 VSS.n2264 0.436245
R9199 VSS.n3549 VSS.n2315 0.436245
R9200 VSS.n3553 VSS.n2316 0.436245
R9201 VSS.n3561 VSS.n2311 0.436245
R9202 VSS.n3566 VSS.n2309 0.436245
R9203 VSS.n5159 VSS.n366 0.436245
R9204 VSS.n5156 VSS.n5155 0.436245
R9205 VSS.n5151 VSS.n374 0.436245
R9206 VSS.n376 VSS.n375 0.436245
R9207 VSS.n3766 VSS.n3757 0.436245
R9208 VSS.n3770 VSS.n3755 0.436245
R9209 VSS.n3775 VSS.n3753 0.436245
R9210 VSS.n3780 VSS.n3751 0.436245
R9211 VSS.n3344 VSS.n3343 0.434398
R9212 VSS.n3208 VSS.n3207 0.434398
R9213 VSS.n3337 VSS.n3213 0.434398
R9214 VSS.n3215 VSS.n3214 0.434398
R9215 VSS.n3325 VSS.n3324 0.434398
R9216 VSS.n3320 VSS.n3227 0.434398
R9217 VSS.n3317 VSS.n3228 0.434398
R9218 VSS.n3314 VSS.n3313 0.434398
R9219 VSS.n3993 VSS.n2120 0.434398
R9220 VSS.n2124 VSS.n2123 0.434398
R9221 VSS.n3988 VSS.n2125 0.434398
R9222 VSS.n3985 VSS.n3984 0.434398
R9223 VSS.n2139 VSS.n2138 0.434398
R9224 VSS.n3975 VSS.n3973 0.434398
R9225 VSS.n2145 VSS.n2144 0.434398
R9226 VSS.n3967 VSS.n2149 0.434398
R9227 VSS.n4597 VSS.n4596 0.434398
R9228 VSS.n1843 VSS.n1842 0.434398
R9229 VSS.n4590 VSS.n1849 0.434398
R9230 VSS.n1851 VSS.n1850 0.434398
R9231 VSS.n4578 VSS.n4577 0.434398
R9232 VSS.n4573 VSS.n1863 0.434398
R9233 VSS.n4570 VSS.n1864 0.434398
R9234 VSS.n4567 VSS.n4566 0.434398
R9235 VSS.n3916 VSS.n2220 0.434398
R9236 VSS.n2353 VSS.n2221 0.434398
R9237 VSS.n2357 VSS.n2351 0.434398
R9238 VSS.n2362 VSS.n2346 0.434398
R9239 VSS.n2371 VSS.n2370 0.434398
R9240 VSS.n2376 VSS.n2375 0.434398
R9241 VSS.n3438 VSS.n2332 0.434398
R9242 VSS.n3436 VSS.n2323 0.434398
R9243 VSS.n4718 VSS.n1622 0.434398
R9244 VSS.n1894 VSS.n1892 0.434398
R9245 VSS.n1941 VSS.n1900 0.434398
R9246 VSS.n1902 VSS.n1901 0.434398
R9247 VSS.n1911 VSS.n1905 0.434398
R9248 VSS.n1927 VSS.n1914 0.434398
R9249 VSS.n1924 VSS.n1919 0.434398
R9250 VSS.n1921 VSS.n1254 0.434398
R9251 VSS.n2535 VSS.n2083 0.433481
R9252 VSS.n2539 VSS.n2533 0.433481
R9253 VSS.n2575 VSS.n2574 0.433481
R9254 VSS.n2570 VSS.n2544 0.433481
R9255 VSS.n2565 VSS.n2551 0.433481
R9256 VSS.n2562 VSS.n2561 0.433481
R9257 VSS.n2557 VSS.n2556 0.433481
R9258 VSS.n3150 VSS.n3147 0.433481
R9259 VSS.n3374 VSS.n3373 0.433481
R9260 VSS.n3369 VSS.n2489 0.433481
R9261 VSS.n3244 VSS.n2491 0.433481
R9262 VSS.n3249 VSS.n3248 0.433481
R9263 VSS.n3258 VSS.n3257 0.433481
R9264 VSS.n3262 VSS.n3261 0.433481
R9265 VSS.n3267 VSS.n3266 0.433481
R9266 VSS.n3382 VSS.n3379 0.433481
R9267 VSS.n3431 VSS.n2396 0.433481
R9268 VSS.n2866 VSS.n2400 0.433481
R9269 VSS.n2871 VSS.n2870 0.433481
R9270 VSS.n2876 VSS.n2875 0.433481
R9271 VSS.n2885 VSS.n2884 0.433481
R9272 VSS.n2889 VSS.n2888 0.433481
R9273 VSS.n2894 VSS.n2893 0.433481
R9274 VSS.n2900 VSS.n2897 0.433481
R9275 VSS.n4627 VSS.n4626 0.433481
R9276 VSS.n4622 VSS.n1827 0.433481
R9277 VSS.n4403 VSS.n1829 0.433481
R9278 VSS.n4408 VSS.n4407 0.433481
R9279 VSS.n4417 VSS.n4416 0.433481
R9280 VSS.n4421 VSS.n4420 0.433481
R9281 VSS.n4426 VSS.n4425 0.433481
R9282 VSS.n4432 VSS.n4429 0.433481
R9283 VSS.n1668 VSS.n1644 0.433481
R9284 VSS.n4713 VSS.n1645 0.433481
R9285 VSS.n1792 VSS.n1790 0.433481
R9286 VSS.n1798 VSS.n1797 0.433481
R9287 VSS.n1809 VSS.n1808 0.433481
R9288 VSS.n1813 VSS.n1812 0.433481
R9289 VSS.n1823 VSS.n1816 0.433481
R9290 VSS.n1821 VSS.n1818 0.433481
R9291 VSS.n5434 VSS.n102 0.433481
R9292 VSS.n5406 VSS.n106 0.433481
R9293 VSS.n133 VSS.n132 0.433481
R9294 VSS.n5401 VSS.n134 0.433481
R9295 VSS.n5393 VSS.n144 0.433481
R9296 VSS.n148 VSS.n147 0.433481
R9297 VSS.n5388 VSS.n149 0.433481
R9298 VSS.n5385 VSS.n5384 0.433481
R9299 VSS.n5141 VSS.n398 0.433481
R9300 VSS.n5113 VSS.n402 0.433481
R9301 VSS.n633 VSS.n632 0.433481
R9302 VSS.n5108 VSS.n634 0.433481
R9303 VSS.n5100 VSS.n644 0.433481
R9304 VSS.n648 VSS.n647 0.433481
R9305 VSS.n5095 VSS.n649 0.433481
R9306 VSS.n5092 VSS.n5091 0.433481
R9307 VSS.n3910 VSS.n3909 0.433481
R9308 VSS.n3905 VSS.n2247 0.433481
R9309 VSS.n3474 VSS.n2249 0.433481
R9310 VSS.n3479 VSS.n3478 0.433481
R9311 VSS.n3493 VSS.n3489 0.433481
R9312 VSS.n3490 VSS.n3467 0.433481
R9313 VSS.n3505 VSS.n3503 0.433481
R9314 VSS.n3510 VSS.n3465 0.433481
R9315 VSS.n4913 VSS.n783 0.433481
R9316 VSS.n4885 VSS.n787 0.433481
R9317 VSS.n840 VSS.n839 0.433481
R9318 VSS.n4880 VSS.n841 0.433481
R9319 VSS.n4872 VSS.n851 0.433481
R9320 VSS.n855 VSS.n854 0.433481
R9321 VSS.n4867 VSS.n856 0.433481
R9322 VSS.n4864 VSS.n4863 0.433481
R9323 VSS.n4772 VSS.n4771 0.433481
R9324 VSS.n4767 VSS.n1280 0.433481
R9325 VSS.n1417 VSS.n1281 0.433481
R9326 VSS.n1422 VSS.n1421 0.433481
R9327 VSS.n1436 VSS.n1412 0.433481
R9328 VSS.n1441 VSS.n1411 0.433481
R9329 VSS.n1444 VSS.n1410 0.433481
R9330 VSS.n1481 VSS.n1449 0.433481
R9331 VSS VSS.n32 0.300074
R9332 VSS VSS.n77 0.300074
R9333 VSS.n3689 VSS 0.300074
R9334 VSS.n1600 VSS 0.300074
R9335 VSS.n1365 VSS 0.300074
R9336 VSS.n1067 VSS 0.300074
R9337 VSS.n4918 VSS 0.300074
R9338 VSS.n3627 VSS 0.300074
R9339 VSS.n3537 VSS 0.300074
R9340 VSS.n5146 VSS 0.300074
R9341 VSS.n3332 VSS 0.298805
R9342 VSS.n2135 VSS 0.298805
R9343 VSS.n4585 VSS 0.298805
R9344 VSS.n2348 VSS 0.298805
R9345 VSS.n1936 VSS 0.298805
R9346 VSS VSS.n2546 0.298174
R9347 VSS VSS.n3252 0.298174
R9348 VSS VSS.n2879 0.298174
R9349 VSS VSS.n4411 0.298174
R9350 VSS VSS.n1801 0.298174
R9351 VSS.n5398 VSS 0.298174
R9352 VSS.n5105 VSS 0.298174
R9353 VSS VSS.n3482 0.298174
R9354 VSS.n4877 VSS 0.298174
R9355 VSS.n1433 VSS 0.298174
R9356 VSS VSS.n0 0.27284
R9357 VSS.n5215 VSS 0.27284
R9358 VSS.n5261 VSS 0.27284
R9359 VSS.n5307 VSS 0.27284
R9360 VSS VSS.n4806 0.27284
R9361 VSS VSS.n4295 0.268748
R9362 VSS VSS.n4315 0.206282
R9363 VSS.n464 VSS 0.13667
R9364 VSS.n545 VSS 0.13667
R9365 VSS.n3694 VSS 0.13667
R9366 VSS.n1311 VSS 0.13667
R9367 VSS VSS.n1364 0.13667
R9368 VSS VSS.n1063 0.13667
R9369 VSS.n1133 VSS 0.13667
R9370 VSS.n2290 VSS 0.13667
R9371 VSS.n3547 VSS 0.13667
R9372 VSS.n3761 VSS 0.13667
R9373 VSS.n3223 VSS 0.136093
R9374 VSS.n3980 VSS 0.136093
R9375 VSS.n1859 VSS 0.136093
R9376 VSS.n2366 VSS 0.136093
R9377 VSS VSS.n1933 0.136093
R9378 VSS.n2547 VSS 0.135807
R9379 VSS.n3253 VSS 0.135807
R9380 VSS.n2880 VSS 0.135807
R9381 VSS.n4412 VSS 0.135807
R9382 VSS.n1803 VSS 0.135807
R9383 VSS VSS.n5397 0.135807
R9384 VSS VSS.n5104 0.135807
R9385 VSS.n3483 VSS 0.135807
R9386 VSS VSS.n4876 0.135807
R9387 VSS VSS.n1432 0.135807
R9388 VSS.n4298 VSS 0.109077
R9389 VSS VSS.n0 0.0549681
R9390 VSS.n5215 VSS 0.0549681
R9391 VSS.n5261 VSS 0.0549681
R9392 VSS.n5307 VSS 0.0549681
R9393 VSS.n4806 VSS 0.0549681
R9394 VSS.n4133 VSS.n4089 0.027734
R9395 VSS.n464 VSS 0.027734
R9396 VSS.n4191 VSS.n4190 0.027734
R9397 VSS.n545 VSS 0.027734
R9398 VSS.n3694 VSS 0.027734
R9399 VSS.n1311 VSS 0.027734
R9400 VSS.n1364 VSS 0.027734
R9401 VSS.n1063 VSS 0.027734
R9402 VSS VSS.n1133 0.027734
R9403 VSS.n2290 VSS 0.027734
R9404 VSS VSS.n3547 0.027734
R9405 VSS VSS.n3761 0.027734
R9406 VSS.n3223 VSS 0.0276186
R9407 VSS.n3980 VSS 0.0276186
R9408 VSS.n1859 VSS 0.0276186
R9409 VSS VSS.n2366 0.0276186
R9410 VSS.n1933 VSS 0.0276186
R9411 VSS.n4271 VSS.n4270 0.0275781
R9412 VSS.n4013 VSS.n4012 0.0275613
R9413 VSS.n2547 VSS 0.0275613
R9414 VSS.n3253 VSS 0.0275613
R9415 VSS.n2880 VSS 0.0275613
R9416 VSS.n4412 VSS 0.0275613
R9417 VSS VSS.n1803 0.0275613
R9418 VSS.n4684 VSS.n4683 0.0275613
R9419 VSS.n4221 VSS.n127 0.0275613
R9420 VSS.n5397 VSS 0.0275613
R9421 VSS.n5104 VSS 0.0275613
R9422 VSS.n3483 VSS 0.0275613
R9423 VSS.n4876 VSS 0.0275613
R9424 VSS.n1432 VSS 0.0275613
R9425 VSS.n1488 VSS.n1487 0.0275613
R9426 VSS.n4272 VSS.n4236 0.0232273
R9427 VSS.n4307 VSS 0.0196718
R9428 VSS.n4246 VSS.n4245 0.00569031
R9429 VSS.n4288 VSS.n4241 0.00134175
R9430 Vbgr.n4 Vbgr.n3 275.454
R9431 Vbgr Vbgr.t0 23.0517
R9432 Vbgr.n5 Vbgr.n4 8.59898
R9433 Vbgr.n0 Vbgr.t3 4.9747
R9434 Vbgr.n2 Vbgr.t6 4.91993
R9435 Vbgr.n1 Vbgr.t5 4.91993
R9436 Vbgr.n0 Vbgr.t4 4.91993
R9437 Vbgr.n3 Vbgr.t2 2.857
R9438 Vbgr.n3 Vbgr.t1 2.857
R9439 Vbgr.n4 Vbgr 2.28652
R9440 Vbgr Vbgr.n2 0.182248
R9441 Vbgr Vbgr.n5 0.0633049
R9442 Vbgr.n5 Vbgr 0.063
R9443 Vbgr.n2 Vbgr.n1 0.0552707
R9444 Vbgr.n1 Vbgr.n0 0.0552707
R9445 MINUS.n6 MINUS.n4 280.998
R9446 MINUS.n1 MINUS.n0 83.5719
R9447 MINUS.n10 MINUS.n9 83.5719
R9448 MINUS.n13 MINUS.n1 73.8498
R9449 MINUS.n5 MINUS.t4 67.4131
R9450 MINUS.n5 MINUS.t5 66.1779
R9451 MINUS.t1 MINUS.n8 64.5544
R9452 MINUS.n9 MINUS.n1 26.074
R9453 MINUS MINUS.n5 11.5195
R9454 MINUS.n6 MINUS.t0 10.2618
R9455 MINUS.n7 MINUS.n6 3.81404
R9456 MINUS.n4 MINUS.t2 2.857
R9457 MINUS.n4 MINUS.t3 2.857
R9458 MINUS.n6 MINUS 2.00868
R9459 MINUS.n12 MINUS.n11 1.5505
R9460 MINUS.n3 MINUS.n2 1.5505
R9461 MINUS.n8 MINUS.n7 1.49631
R9462 MINUS.n8 MINUS.n3 1.41981
R9463 MINUS.n10 MINUS.n3 1.07024
R9464 MINUS.n11 MINUS.n0 0.885803
R9465 MINUS.n11 MINUS.n10 0.77514
R9466 MINUS MINUS.n0 0.756696
R9467 MINUS.n13 MINUS.n12 0.71401
R9468 MINUS MINUS.n13 0.576402
R9469 MINUS.n9 MINUS.t1 0.290206
R9470 MINUS.n12 MINUS.n2 0.0205321
R9471 MINUS.n7 MINUS.n2 0.00130128
R9472 Gcm1.n0 Gcm1.t4 289.291
R9473 Gcm1.n0 Gcm1.t0 288.884
R9474 Gcm1.n2 Gcm1.t1 231.746
R9475 Gcm1.n2 Gcm1.n1 211.613
R9476 Gcm1 Gcm1.n2 5.53507
R9477 Gcm1 Gcm1.n0 5.21741
R9478 Gcm1.n1 Gcm1.t3 2.1755
R9479 Gcm1.n1 Gcm1.t2 2.1755
C0 a_23884_n8277# a_24050_n8277# 0.432514f
C1 a_24216_n8877# a_25472_n8877# 0.001551f
C2 Vbgr a_24605_n9724# 1.13e-19
C3 Gcm1 MINUS 0.027313f
C4 XQ2[0|0].Emitter a_25307_n10376# 0.003384f
C5 Sop Gcm2 0.109242f
C6 a_24137_n9724# a_24371_n10376# 0.034612f
C7 a_24050_n8277# Gcm2 8.48e-19
C8 a_24808_n8877# PLUS 0.003696f
C9 XQ2[0|0].Emitter VDD 0.264478f
C10 a_23552_n8877# XQ2[0|0].Emitter 0.004761f
C11 a_24808_n8877# a_24974_n8277# 0.023915f
C12 Sop PLUS 1.98461f
C13 Vbgr a_25307_n10376# 0.033913f
C14 a_23669_n9724# a_23552_n8877# 0.042257f
C15 a_23884_n8277# XQ2[0|0].Emitter 0.001537f
C16 a_23718_n8877# XQ2[0|0].Emitter 0.002687f
C17 a_24050_n8277# PLUS 0.118024f
C18 a_24808_n8877# MINUS 0.005358f
C19 XQ2[0|0].Emitter Vbgr 0.766448f
C20 a_23884_n8277# VDD 3.52e-19
C21 a_24839_n10376# a_24371_n10376# 0.298765f
C22 a_25307_n10376# a_23903_n10376# 1.89e-21
C23 a_23552_n8877# a_23884_n8277# 0.003644f
C24 VDD Vbgr 3.58636f
C25 a_23552_n8877# a_23718_n8877# 0.745688f
C26 a_24371_n10376# a_24605_n9724# 0.034601f
C27 a_24216_n8877# a_24137_n9724# 0.033727f
C28 Sop MINUS 1.89228f
C29 a_23669_n9724# Vbgr 3.15e-21
C30 Gcm2 XQ2[0|0].Emitter 0.024343f
C31 a_24839_n10376# a_25073_n9724# 0.034607f
C32 Gcm2 VDD 1.05773f
C33 a_24050_n8277# MINUS 0.004852f
C34 a_23552_n8877# a_23903_n10376# 0.003748f
C35 a_25073_n9724# a_24605_n9724# 0.29801f
C36 a_24216_n8877# a_24808_n8877# 0.453352f
C37 a_23552_n8877# Gcm2 0.002655f
C38 a_23718_n8877# a_23884_n8277# 0.023433f
C39 a_23669_n9724# a_23903_n10376# 0.034605f
C40 a_23669_n9724# Gcm2 4.78e-20
C41 PLUS XQ2[0|0].Emitter 0.041558f
C42 a_25307_n10376# a_24371_n10376# 4.82e-21
C43 a_23884_n8277# Gcm2 0.055631f
C44 a_24216_n8877# a_24839_n10376# 0.004947f
C45 a_23718_n8877# Gcm2 0.004231f
C46 a_24974_n8277# XQ2[0|0].Emitter 9.61e-19
C47 PLUS VDD 1.05274f
C48 Gcm2 Vbgr 0.005993f
C49 a_24216_n8877# a_24605_n9724# 0.042461f
C50 a_24050_n8277# a_24216_n8877# 0.023433f
C51 XQ2[0|0].Emitter a_24371_n10376# 0.002121f
C52 MINUS a_25307_n10376# 1.23e-19
C53 a_25073_n9724# a_25307_n10376# 0.034603f
C54 a_23435_n10376# a_24839_n10376# 3.11e-21
C55 MINUS XQ2[0|0].Emitter 4.74122f
C56 a_25140_n8277# XQ2[0|0].Emitter 9.32e-19
C57 XQ2[0|0].Emitter a_25073_n9724# 0.058405f
C58 a_23884_n8277# PLUS 0.317764f
C59 a_23718_n8877# PLUS 1.02e-20
C60 MINUS VDD 0.940915f
C61 PLUS Vbgr 0.058292f
C62 a_23552_n8877# MINUS 0.001132f
C63 a_23884_n8277# a_24974_n8277# 0.340116f
C64 Sop Gcm1 0.18188f
C65 Gcm2 PLUS 1.2386f
C66 a_24216_n8877# XQ2[0|0].Emitter 0.381626f
C67 a_23884_n8277# MINUS 0.026861f
C68 a_23718_n8877# MINUS 0.001041f
C69 a_23386_n8277# a_23552_n8877# 0.023433f
C70 a_23903_n10376# a_24371_n10376# 0.298666f
C71 a_25472_n8877# a_25307_n10376# 0.002985f
C72 MINUS Vbgr 0.428769f
C73 Vbgr a_25073_n9724# 0.297712f
C74 a_23435_n10376# a_25307_n10376# 6.09e-22
C75 a_23552_n8877# a_24216_n8877# 0.337637f
C76 a_25472_n8877# XQ2[0|0].Emitter 0.017877f
C77 Gcm2 MINUS 0.65619f
C78 a_23386_n8277# a_23884_n8277# 1.41e-19
C79 a_24137_n9724# a_24605_n9724# 0.298808f
C80 a_24050_n8277# a_24137_n9724# 0.002284f
C81 a_23386_n8277# Vbgr 2.71e-19
C82 a_23435_n10376# a_23552_n8877# 0.004809f
C83 a_23884_n8277# a_24216_n8877# 0.017118f
C84 a_24974_n8277# PLUS 0.499589f
C85 a_23435_n10376# a_23669_n9724# 0.034723f
C86 a_24216_n8877# Vbgr 2.61e-19
C87 a_23386_n8277# Gcm2 0.021107f
C88 PLUS MINUS 2.82036f
C89 a_25472_n8877# Vbgr 0.030096f
C90 a_24216_n8877# Gcm2 4.84e-19
C91 a_25140_n8277# PLUS 0.002742f
C92 Gcm1 VDD 2.09957f
C93 a_24974_n8277# MINUS 0.213061f
C94 a_24974_n8277# a_25140_n8277# 0.737085f
C95 a_24974_n8277# a_25073_n9724# 0.001698f
C96 a_24839_n10376# a_24605_n9724# 0.034601f
C97 a_23435_n10376# a_23903_n10376# 0.298736f
C98 a_23386_n8277# PLUS 0.001339f
C99 a_24216_n8877# PLUS 1.75e-19
C100 a_25140_n8277# MINUS 0.068246f
C101 MINUS a_25073_n9724# 0.00849f
C102 Gcm1 Vbgr 4.69e-19
C103 a_25140_n8277# a_25073_n9724# 0.003106f
C104 a_24216_n8877# a_24974_n8277# 0.003676f
C105 a_23669_n9724# a_24137_n9724# 0.298213f
C106 a_24808_n8877# XQ2[0|0].Emitter 0.112162f
C107 a_24216_n8877# a_24371_n10376# 0.004861f
C108 a_25472_n8877# PLUS 0.025645f
C109 a_23386_n8277# MINUS 0.006469f
C110 a_24974_n8277# a_25472_n8877# 0.023915f
C111 a_24839_n10376# a_25307_n10376# 0.299281f
C112 a_24216_n8877# MINUS 0.349768f
C113 a_24216_n8877# a_25140_n8277# 0.023915f
C114 a_24216_n8877# a_25073_n9724# 0.015496f
C115 Vbgr a_24137_n9724# 1.56e-20
C116 a_23435_n10376# a_24371_n10376# 7.87e-20
C117 XQ2[0|0].Emitter a_24839_n10376# 0.003391f
C118 Sop VDD 9.75e-19
C119 XQ2[0|0].Emitter a_24605_n9724# 0.059011f
C120 a_25472_n8877# MINUS 0.514607f
C121 a_23884_n8277# a_24808_n8877# 0.023915f
C122 a_23903_n10376# a_24137_n9724# 0.034611f
C123 Gcm1 PLUS 0.4684f
C124 Gcm2 a_24137_n9724# 1.86e-20
C125 a_23552_n8877# a_24050_n8277# 0.023451f
C126 Vbgr VSS 13.494073f
C127 VDD VSS 33.08502f
C128 a_25307_n10376# VSS 0.806369f
C129 a_25073_n9724# VSS 0.467234f
C130 a_24839_n10376# VSS 0.505692f
C131 a_24605_n9724# VSS 0.462354f
C132 a_24371_n10376# VSS 0.505614f
C133 a_24137_n9724# VSS 0.466284f
C134 a_23903_n10376# VSS 0.506957f
C135 a_23669_n9724# VSS 0.754256f
C136 a_23435_n10376# VSS 0.837674f
C137 a_25472_n8877# VSS 0.640408f
C138 a_25140_n8277# VSS 0.315247f
C139 a_24974_n8277# VSS 0.437807f
C140 a_24808_n8877# VSS 0.472164f
C141 a_24216_n8877# VSS 0.820643f
C142 a_24050_n8277# VSS 0.450227f
C143 a_23884_n8277# VSS 1.14965f
C144 a_23718_n8877# VSS 0.336042f
C145 a_23552_n8877# VSS 0.815395f
C146 a_23386_n8277# VSS 0.987226f
C147 Sop VSS 2.73918f
C148 XQ2[0|0].Emitter VSS 77.905106f
C149 MINUS VSS 7.324422f
C150 PLUS VSS 7.04395f
C151 Gcm2 VSS 5.54568f
C152 Gcm1 VSS 2.196767f
C153 Gcm1.t4 VSS 0.399998f
C154 Gcm1.t0 VSS 0.39981f
C155 Gcm1.n0 VSS 0.271096f
C156 Gcm1.t3 VSS 0.034704f
C157 Gcm1.t2 VSS 0.034704f
C158 Gcm1.n1 VSS 0.123204f
C159 Gcm1.t1 VSS 0.185044f
C160 Gcm1.n2 VSS 0.445974f
C161 MINUS.n0 VSS 0.036563f
C162 MINUS.n1 VSS 0.165732f
C163 MINUS.n2 VSS 0.038416f
C164 MINUS.n3 VSS 0.068317f
C165 MINUS.t2 VSS 0.034333f
C166 MINUS.t3 VSS 0.034333f
C167 MINUS.n4 VSS 0.12246f
C168 MINUS.t4 VSS 1.24342f
C169 MINUS.t5 VSS 1.23503f
C170 MINUS.n5 VSS 1.09001f
C171 MINUS.t0 VSS 0.113521f
C172 MINUS.n6 VSS 0.940622f
C173 MINUS.n7 VSS 0.876222f
C174 MINUS.n8 VSS 0.193729f
C175 MINUS.t1 VSS 0.135718f
C176 MINUS.n9 VSS 0.03663f
C177 MINUS.n10 VSS 0.041082f
C178 MINUS.n11 VSS 0.036974f
C179 MINUS.n12 VSS 0.274275f
C180 MINUS.n13 VSS 0.187128f
C181 Vbgr.t3 VSS 0.998618f
C182 Vbgr.t4 VSS 0.985768f
C183 Vbgr.n0 VSS 2.36767f
C184 Vbgr.t5 VSS 0.985768f
C185 Vbgr.n1 VSS 1.21061f
C186 Vbgr.t6 VSS 0.985768f
C187 Vbgr.n2 VSS 1.17183f
C188 Vbgr.t0 VSS 0.058596f
C189 Vbgr.t2 VSS 0.046655f
C190 Vbgr.t1 VSS 0.046655f
C191 Vbgr.n3 VSS 0.161469f
C192 Vbgr.n4 VSS 0.897488f
C193 Vbgr.n5 VSS 0.835527f
C194 VDD.n0 VSS 0.101411f
C195 VDD.n1 VSS 0.192556f
C196 VDD.t6 VSS 0.125212f
C197 VDD.n2 VSS 0.100291f
C198 VDD.t2 VSS 0.125172f
C199 VDD.t8 VSS 0.141798f
C200 VDD.t18 VSS 0.022103f
C201 VDD.n3 VSS 0.076481f
C202 VDD.n4 VSS 0.093741f
C203 VDD.t10 VSS 0.022103f
C204 VDD.t14 VSS 0.022103f
C205 VDD.n5 VSS 0.076481f
C206 VDD.n6 VSS 0.087797f
C207 VDD.t20 VSS 0.022103f
C208 VDD.t24 VSS 0.022103f
C209 VDD.n7 VSS 0.076481f
C210 VDD.n8 VSS 0.087797f
C211 VDD.t12 VSS 0.022103f
C212 VDD.t16 VSS 0.022103f
C213 VDD.n9 VSS 0.076481f
C214 VDD.n10 VSS 0.087797f
C215 VDD.t22 VSS 0.022103f
C216 VDD.t4 VSS 0.022103f
C217 VDD.n11 VSS 0.076481f
C218 VDD.n12 VSS 0.094769f
C219 VDD.n13 VSS 0.101331f
C220 VDD.n14 VSS 0.048367f
C221 VDD.t5 VSS 0.119696f
C222 VDD.n15 VSS 0.194388f
C223 VDD.n16 VSS 0.483776f
C224 VDD.t3 VSS 0.430292f
C225 VDD.t21 VSS 0.260354f
C226 VDD.t15 VSS 0.260354f
C227 VDD.t11 VSS 0.260354f
C228 VDD.t23 VSS 0.260354f
C229 VDD.t19 VSS 0.260354f
C230 VDD.t13 VSS 0.260354f
C231 VDD.t9 VSS 0.260354f
C232 VDD.t17 VSS 0.260354f
C233 VDD.t7 VSS 0.407816f
C234 VDD.n17 VSS 0.321909f
C235 VDD.n18 VSS 0.049622f
C236 VDD.n19 VSS 0.213927f
C237 VDD.n20 VSS 0.440923f
C238 VDD.t25 VSS 0.674994f
C239 VDD.t0 VSS 0.660024f
C240 VDD.n21 VSS 0.701578f
C241 VDD.t26 VSS 0.017682f
C242 VDD.t1 VSS 0.017682f
C243 VDD.n22 VSS 0.060101f
C244 VDD.n23 VSS 0.185965f
C245 VDD.n24 VSS 0.810651f
C246 VDD.n25 VSS 0.125027f
C247 VDD.n26 VSS 0.261933f
C248 PLUS.t2 VSS 0.019129f
C249 PLUS.t3 VSS 0.019129f
C250 PLUS.n0 VSS 0.066396f
C251 PLUS.t1 VSS 0.020814f
C252 PLUS.t0 VSS 0.008975f
C253 PLUS.n1 VSS 0.195549f
C254 PLUS.n2 VSS 0.201296f
C255 PLUS.t5 VSS 0.692798f
C256 PLUS.t4 VSS 0.688119f
C257 PLUS.n3 VSS 0.530095f
C258 opout.n0 VSS 1.7936f
C259 opout.n1 VSS 1.60492f
C260 opout.t6 VSS 0.015326f
C261 opout.t2 VSS 0.015129f
C262 opout.t5 VSS 1.82387f
C263 opout.t1 VSS 1.11063f
C264 opout.t3 VSS 1.82387f
C265 opout.t7 VSS 1.11063f
C266 opout.n2 VSS 0.969049f
C267 opout.t8 VSS 0.015129f
C268 opout.t4 VSS 0.015129f
C269 opout.t14 VSS 0.233109f
C270 opout.t18 VSS 0.233099f
C271 opout.t16 VSS 0.233099f
C272 opout.t13 VSS 0.233099f
C273 opout.t11 VSS 0.233099f
C274 opout.t17 VSS 0.233099f
C275 opout.t15 VSS 0.233099f
C276 opout.t12 VSS 0.233099f
C277 opout.t0 VSS 0.032942f
C278 opout.t9 VSS 0.032942f
C279 opout.n3 VSS 0.116455f
C280 opout.t10 VSS 0.176215f
C281 opout.n4 VSS 0.479365f
.ends

