magic
tech sky130A
magscale 1 2
timestamp 1725582067
<< nwell >>
rect 7885 -7401 8086 -7396
rect 7885 -9194 10486 -7401
rect 18117 -8602 21539 -8594
rect 8081 -9204 10486 -9194
rect 17995 -10396 21799 -8602
rect 17995 -10404 18211 -10396
rect 18631 -13251 20855 -12387
rect 18619 -15729 20843 -15717
rect 18619 -16127 18637 -15729
rect 20825 -16127 20843 -15729
rect 18619 -16593 20843 -16127
<< pwell >>
rect 12395 -5817 12660 -5625
rect 12589 -5824 12659 -5817
rect 12918 -5834 12993 -5466
rect 13416 -5818 13489 -5446
rect 12918 -6779 12993 -6411
rect 13253 -6774 13324 -6425
rect 13748 -6774 13819 -6427
rect 13910 -6779 13985 -6411
rect 14572 -6625 14845 -6395
rect 12515 -9868 12731 -9404
rect 12515 -10469 12731 -10005
rect 12987 -10493 13203 -10029
rect 18373 -10967 18743 -10965
rect 18211 -11394 18743 -10967
<< nbase >>
rect 12716 -13745 12717 -13706
<< pmoslvt >>
rect 18743 -13139 20743 -12939
<< pdiff >>
rect 18685 -12951 18743 -12939
rect 18685 -13127 18697 -12951
rect 18731 -13127 18743 -12951
rect 18685 -13139 18743 -13127
rect 20743 -12951 20801 -12939
rect 20743 -13127 20755 -12951
rect 20789 -13127 20801 -12951
rect 20743 -13139 20801 -13127
rect 12716 -13745 12717 -13706
<< pdiffc >>
rect 18697 -13127 18731 -12951
rect 20755 -13127 20789 -12951
<< psubdiff >>
rect 22996 -3003 23983 -2979
rect 6004 -3990 6028 -3003
rect 23983 -3990 24007 -3003
rect 10684 -7265 10880 -7208
rect 10684 -8547 10732 -7265
rect 10846 -8547 10880 -7265
rect 10684 -8605 10880 -8547
rect 16490 -7258 16686 -7201
rect 16490 -8540 16538 -7258
rect 16652 -8540 16686 -7258
rect 16490 -8598 16686 -8540
rect 17811 -8189 17931 -8104
rect 17811 -8689 17851 -8189
rect 17896 -8689 17931 -8189
rect 17811 -8799 17931 -8689
rect 6004 -18983 6028 -17996
rect 23983 -18983 24007 -17996
rect 22996 -19007 23983 -18983
<< nsubdiff >>
rect 8030 -7877 8240 -7803
rect 8030 -8737 8076 -7877
rect 8170 -8737 8240 -7877
rect 8030 -8802 8240 -8737
rect 10141 -7867 10351 -7793
rect 10141 -8727 10187 -7867
rect 10281 -8727 10351 -7867
rect 10141 -8792 10351 -8727
rect 18066 -9091 18262 -9030
rect 18066 -10148 18114 -9091
rect 18201 -10148 18262 -9091
rect 18066 -10202 18262 -10148
rect 21426 -9071 21622 -9010
rect 21426 -10128 21474 -9071
rect 21561 -10128 21622 -9071
rect 21426 -10182 21622 -10128
rect 18891 -12570 20642 -12509
rect 18891 -12669 19075 -12570
rect 20472 -12669 20642 -12570
rect 18891 -12730 20642 -12669
rect 18832 -16311 20583 -16250
rect 18832 -16410 19002 -16311
rect 20399 -16410 20583 -16311
rect 18832 -16471 20583 -16410
<< psubdiffcont >>
rect 6028 -3990 23983 -3003
rect 6028 -17996 7015 -3990
rect 10732 -8547 10846 -7265
rect 16538 -8540 16652 -7258
rect 17851 -8689 17896 -8189
rect 22996 -17996 23983 -3990
rect 6028 -18983 23983 -17996
<< nsubdiffcont >>
rect 8076 -8737 8170 -7877
rect 10187 -8727 10281 -7867
rect 18114 -10148 18201 -9091
rect 21474 -10128 21561 -9071
rect 19075 -12669 20472 -12570
rect 19002 -16410 20399 -16311
<< poly >>
rect 18743 -12858 20743 -12842
rect 18743 -12892 18759 -12858
rect 20727 -12892 20743 -12858
rect 18743 -12939 20743 -12892
rect 18743 -13186 20743 -13139
rect 18743 -13220 18759 -13186
rect 20727 -13220 20743 -13186
rect 18743 -13236 20743 -13220
<< polycont >>
rect 18759 -12892 20727 -12858
rect 18759 -13220 20727 -13186
<< locali >>
rect 22996 -3003 23983 -2987
rect 6012 -3990 6028 -3003
rect 23983 -3990 23999 -3003
rect 10710 -7265 10863 -7237
rect 8058 -7877 8193 -7840
rect 8058 -7943 8076 -7877
rect 8170 -7943 8193 -7877
rect 10169 -7867 10304 -7830
rect 10169 -7941 10187 -7867
rect 10281 -7941 10304 -7867
rect 8192 -8200 8193 -7943
rect 10710 -8188 10716 -7265
rect 8058 -8737 8076 -8200
rect 8170 -8737 8193 -8200
rect 8058 -8760 8193 -8737
rect 10169 -8727 10187 -8200
rect 10281 -8727 10304 -8200
rect 10846 -8188 10863 -7265
rect 16516 -7258 16669 -7230
rect 16516 -7265 16538 -7258
rect 16652 -7265 16669 -7258
rect 16516 -8214 16537 -7265
rect 16667 -8214 16669 -7265
rect 17831 -8189 17901 -8149
rect 17831 -8299 17851 -8189
rect 17896 -8299 17901 -8189
rect 16516 -8568 16669 -8566
rect 17831 -8689 17851 -8499
rect 17896 -8689 17901 -8499
rect 17831 -8724 17901 -8689
rect 10169 -8750 10304 -8727
rect 18226 -9331 18228 -9064
rect 18100 -10148 18114 -9331
rect 18201 -10148 18228 -9331
rect 21460 -10128 21474 -9335
rect 21561 -10128 21588 -9335
rect 21460 -10148 21588 -10128
rect 18100 -10168 18228 -10148
rect 9809 -17137 10044 -10766
rect 9826 -17196 10044 -17137
rect 10862 -16791 11276 -10757
rect 12216 -10762 12506 -10756
rect 12216 -10841 13214 -10762
rect 13379 -10786 14010 -10773
rect 13379 -10840 13973 -10786
rect 10862 -17203 11332 -16791
rect 12216 -16800 12620 -10841
rect 12716 -13745 12717 -13706
rect 10862 -17204 11276 -17203
rect 12147 -17204 12620 -16800
rect 13436 -17203 13909 -10840
rect 14724 -17204 15195 -10761
rect 16012 -17202 16485 -10762
rect 17301 -17137 17537 -10761
rect 18962 -12570 19432 -12556
rect 20063 -12570 20543 -12556
rect 18962 -12669 19075 -12570
rect 20472 -12669 20543 -12570
rect 18962 -12679 19432 -12669
rect 20063 -12679 20543 -12669
rect 18962 -12688 20543 -12679
rect 18743 -12892 18759 -12858
rect 20727 -12892 20743 -12858
rect 18697 -12951 18731 -12935
rect 18697 -13143 18731 -13127
rect 20755 -12951 20789 -12935
rect 20755 -13143 20789 -13127
rect 18743 -13220 18759 -13186
rect 20727 -13220 20743 -13186
rect 18931 -16301 20512 -16292
rect 18931 -16311 19411 -16301
rect 20042 -16311 20512 -16301
rect 18931 -16410 19002 -16311
rect 20399 -16410 20512 -16311
rect 18931 -16424 19411 -16410
rect 20042 -16424 20512 -16410
rect 17301 -17201 17520 -17137
rect 6012 -18983 6028 -17996
rect 23983 -18983 23999 -17996
rect 22996 -18999 23983 -18983
<< viali >>
rect 10637 -3889 10961 -3194
rect 12234 -3866 12419 -3102
rect 14781 -3820 15105 -3125
rect 16309 -3935 16865 -3102
rect 17692 -3629 17735 -3586
rect 12288 -6602 12344 -5605
rect 14892 -6623 14948 -5626
rect 8056 -8200 8076 -7943
rect 8076 -8200 8170 -7943
rect 8170 -8200 8192 -7943
rect 10168 -8200 10187 -7941
rect 10187 -8200 10281 -7941
rect 10281 -8200 10304 -7941
rect 10716 -8188 10732 -7265
rect 10708 -8547 10732 -8188
rect 10732 -8547 10846 -7265
rect 10846 -8547 10865 -8188
rect 16537 -8214 16538 -7265
rect 10708 -8580 10865 -8547
rect 16515 -8540 16538 -8214
rect 16538 -8540 16652 -7265
rect 16652 -8214 16667 -7265
rect 16652 -8540 16669 -8214
rect 17826 -8499 17851 -8299
rect 17851 -8499 17896 -8299
rect 17896 -8499 17911 -8299
rect 16515 -8566 16669 -8540
rect 18096 -9091 18226 -9060
rect 18096 -9331 18114 -9091
rect 18114 -9331 18201 -9091
rect 18201 -9331 18226 -9091
rect 12519 -10472 12587 -9474
rect 13132 -10477 13200 -9478
rect 21453 -9071 21591 -9042
rect 21453 -9335 21474 -9071
rect 21474 -9335 21561 -9071
rect 21561 -9335 21591 -9071
rect 18214 -11383 18282 -10967
rect 21148 -11371 21206 -10966
rect 18214 -12031 18272 -11613
rect 21160 -12016 21218 -11611
rect 19432 -12570 20063 -12533
rect 19432 -12669 20063 -12570
rect 19432 -12679 20063 -12669
rect 19251 -12892 20235 -12858
rect 18697 -13127 18731 -12951
rect 20755 -13127 20789 -12951
rect 19251 -13220 20235 -13186
rect 20883 -14582 20940 -14091
rect 19411 -16311 20042 -16301
rect 19411 -16410 20042 -16311
rect 19411 -16447 20042 -16410
rect 18039 -18727 18385 -18071
<< metal1 >>
rect 12228 -3102 12425 -3090
rect 10631 -3194 10967 -3182
rect 10631 -3889 10637 -3194
rect 10961 -3889 10967 -3194
rect 12228 -3866 12234 -3102
rect 12419 -3866 12425 -3102
rect 16303 -3102 16871 -3090
rect 14775 -3125 15111 -3113
rect 14775 -3820 14781 -3125
rect 15105 -3820 15111 -3125
rect 14775 -3832 15111 -3820
rect 12228 -3878 12425 -3866
rect 10631 -3901 10967 -3889
rect 10683 -7265 10868 -3901
rect 12280 -5605 12350 -3878
rect 12920 -5466 13325 -5449
rect 12280 -6602 12288 -5605
rect 12344 -5626 12350 -5605
rect 12918 -5524 13325 -5466
rect 12395 -5626 12660 -5625
rect 12344 -5817 12660 -5626
rect 12344 -6015 12500 -5817
rect 12589 -5824 12659 -5817
rect 12741 -5827 12751 -5607
rect 12822 -5827 12832 -5607
rect 12918 -5834 12993 -5524
rect 13075 -5829 13085 -5609
rect 13156 -5829 13166 -5609
rect 13250 -5817 13325 -5524
rect 13416 -5519 13986 -5446
rect 13416 -5818 13489 -5519
rect 13737 -5831 13747 -5611
rect 13818 -5831 13828 -5611
rect 13913 -5825 13986 -5519
rect 14243 -5528 14647 -5453
rect 14070 -5832 14080 -5612
rect 14151 -5832 14161 -5612
rect 14243 -5821 14318 -5528
rect 14399 -5927 14409 -5618
rect 14481 -5927 14491 -5618
rect 14571 -5825 14646 -5528
rect 14897 -5614 14967 -3832
rect 16303 -3935 16309 -3102
rect 16865 -3935 16871 -3102
rect 16303 -3947 16871 -3935
rect 17686 -3586 17741 -3574
rect 17686 -3629 17692 -3586
rect 17735 -3629 17741 -3586
rect 14886 -5619 14967 -5614
rect 14750 -5626 14967 -5619
rect 14750 -6008 14892 -5626
rect 12344 -6234 12350 -6015
rect 12344 -6602 12493 -6234
rect 12280 -6621 12493 -6602
rect 12295 -6623 12493 -6621
rect 12585 -6700 12660 -6411
rect 12741 -6648 12751 -6212
rect 12829 -6648 12839 -6212
rect 14886 -6234 14892 -6008
rect 14750 -6395 14892 -6234
rect 12918 -6700 12993 -6411
rect 13075 -6643 13085 -6423
rect 13156 -6643 13166 -6423
rect 12585 -6775 12993 -6700
rect 13253 -6702 13324 -6425
rect 13409 -6644 13419 -6424
rect 13490 -6644 13500 -6424
rect 13748 -6702 13819 -6427
rect 13253 -6773 13819 -6702
rect 13910 -6708 13985 -6411
rect 14071 -6645 14081 -6425
rect 14152 -6645 14162 -6425
rect 14243 -6708 14318 -6406
rect 14403 -6645 14413 -6425
rect 14484 -6645 14494 -6425
rect 14572 -6623 14892 -6395
rect 14948 -6623 14967 -5626
rect 14572 -6625 14845 -6623
rect 14886 -6635 14967 -6623
rect 14897 -6667 14967 -6635
rect 13253 -6774 13324 -6773
rect 13748 -6774 13819 -6773
rect 12585 -6779 12660 -6775
rect 12918 -6779 12993 -6775
rect 13909 -6783 14318 -6708
rect 11885 -7119 15489 -7110
rect 8721 -7804 9701 -7798
rect 8050 -7943 8198 -7931
rect 8421 -7943 8651 -7842
rect 8721 -7882 9162 -7804
rect 9152 -7899 9162 -7882
rect 9256 -7882 9701 -7804
rect 9256 -7899 9266 -7882
rect 9763 -7943 10013 -7826
rect 10162 -7941 10310 -7929
rect 10158 -7943 10168 -7941
rect 8046 -8200 8056 -7943
rect 8192 -8200 10168 -7943
rect 10304 -8200 10314 -7941
rect 10683 -8188 10716 -7265
rect 10846 -8176 10868 -7265
rect 11077 -7196 16269 -7119
rect 16342 -7196 16464 -7190
rect 11077 -7318 16342 -7196
rect 11077 -7616 16269 -7318
rect 16342 -7324 16464 -7318
rect 16494 -7265 16679 -3947
rect 10846 -8188 10871 -8176
rect 8050 -8212 8198 -8200
rect 10162 -8212 10310 -8200
rect 10683 -8311 10708 -8188
rect 8651 -8830 8735 -8442
rect 9165 -8707 9175 -8453
rect 9245 -8707 9255 -8453
rect 9683 -8830 9767 -8438
rect 10702 -8580 10708 -8311
rect 10865 -8190 10871 -8188
rect 10865 -8580 11137 -8190
rect 14494 -8272 14500 -8188
rect 14584 -8272 14590 -8188
rect 16494 -8213 16537 -7265
rect 16237 -8214 16537 -8213
rect 16667 -8214 16679 -7265
rect 16801 -7318 16807 -7196
rect 16929 -7318 17285 -7196
rect 12773 -8562 12783 -8289
rect 12847 -8562 12857 -8289
rect 10702 -8592 11137 -8580
rect 10708 -8701 11137 -8592
rect 16237 -8566 16515 -8214
rect 16669 -8332 16679 -8214
rect 16669 -8463 16995 -8332
rect 16669 -8566 16675 -8463
rect 16237 -8578 16675 -8566
rect 16864 -8556 16995 -8463
rect 17163 -8466 17285 -7318
rect 17686 -8319 17741 -3629
rect 17820 -8299 17917 -8287
rect 17820 -8319 17826 -8299
rect 17508 -8462 17518 -8335
rect 17574 -8462 17584 -8335
rect 17686 -8499 17826 -8319
rect 17911 -8499 17917 -8299
rect 17686 -8504 17917 -8499
rect 17686 -8556 17741 -8504
rect 17820 -8511 17917 -8504
rect 10706 -8790 11931 -8701
rect 10706 -8808 10708 -8790
rect 8651 -8914 9767 -8830
rect 9683 -9116 9767 -8914
rect 10936 -8808 11931 -8790
rect 11995 -8816 13647 -8720
rect 11995 -9012 12808 -8816
rect 12968 -9012 13647 -8816
rect 13713 -8810 15365 -8720
rect 16237 -8724 16666 -8578
rect 16864 -8681 17741 -8556
rect 15443 -8763 16668 -8724
rect 15441 -8809 16668 -8763
rect 16864 -8802 16995 -8681
rect 17586 -8714 17741 -8681
rect 17365 -8736 17417 -8730
rect 17097 -8788 17365 -8738
rect 17417 -8743 17519 -8738
rect 17417 -8788 17521 -8743
rect 13713 -9011 14206 -8810
rect 14407 -9011 15365 -8810
rect 15443 -8831 16668 -8809
rect 17097 -8810 17521 -8788
rect 17586 -8795 17734 -8714
rect 13713 -9012 15365 -9011
rect 10708 -9024 10936 -9018
rect 12800 -9017 12808 -9012
rect 12908 -9017 12970 -9012
rect 14117 -9014 14201 -9012
rect 12800 -9024 12970 -9017
rect 9683 -9200 14500 -9116
rect 14584 -9200 14590 -9116
rect 12515 -9415 12731 -9404
rect 12238 -9429 12466 -9423
rect 12513 -9429 12731 -9415
rect 13126 -9428 13206 -9420
rect 12466 -9474 12731 -9429
rect 12466 -9657 12519 -9474
rect 12238 -9663 12466 -9657
rect 12513 -10472 12519 -9657
rect 12587 -9868 12731 -9474
rect 12971 -9478 13206 -9428
rect 12802 -9734 12808 -9634
rect 12908 -9734 12914 -9634
rect 12587 -10005 12593 -9868
rect 12971 -9892 13132 -9478
rect 12587 -10469 12731 -10005
rect 13126 -10029 13132 -9892
rect 12801 -10469 12811 -10157
rect 12899 -10469 12909 -10157
rect 12587 -10472 12593 -10469
rect 12513 -10484 12593 -10472
rect 12987 -10477 13132 -10029
rect 13200 -10477 13206 -9478
rect 17425 -9879 17521 -8810
rect 18580 -8838 21055 -8820
rect 18580 -8892 18832 -8838
rect 20522 -8892 21055 -8838
rect 18368 -9003 18513 -8920
rect 18580 -8979 21055 -8892
rect 21212 -8917 21271 -8915
rect 21128 -8986 21271 -8917
rect 18070 -9044 18273 -9042
rect 18368 -9044 18426 -9003
rect 21212 -9044 21271 -8986
rect 21447 -9042 21597 -9030
rect 21443 -9044 21453 -9042
rect 18070 -9060 21453 -9044
rect 18070 -9331 18096 -9060
rect 18226 -9331 21453 -9060
rect 18090 -9333 21453 -9331
rect 18090 -9343 18232 -9333
rect 17425 -9975 17980 -9879
rect 13427 -10169 13433 -9994
rect 13608 -10169 17135 -9994
rect 17310 -10169 17316 -9994
rect 12987 -10489 13206 -10477
rect 17884 -10431 17980 -9975
rect 18368 -9997 18426 -9333
rect 19753 -9487 21116 -9480
rect 19753 -9591 21142 -9487
rect 18666 -10342 18760 -9677
rect 18982 -9988 19070 -9677
rect 19285 -9796 19295 -9650
rect 19405 -9796 19415 -9650
rect 19759 -9663 19870 -9591
rect 19629 -9671 20019 -9663
rect 19303 -9822 19393 -9796
rect 18909 -9994 19084 -9988
rect 18909 -10175 19084 -10169
rect 19303 -10145 19391 -9822
rect 19621 -9990 20019 -9671
rect 20230 -9792 20240 -9659
rect 20359 -9792 20369 -9659
rect 19623 -10022 20019 -9990
rect 19629 -10027 20019 -10022
rect 20251 -10145 20339 -9792
rect 20561 -9988 20649 -9680
rect 18668 -10431 18760 -10342
rect 18982 -10313 19070 -10175
rect 19303 -10233 20339 -10145
rect 20494 -9994 20669 -9988
rect 20494 -10175 20669 -10169
rect 20561 -10313 20649 -10175
rect 18982 -10401 20649 -10313
rect 20881 -10431 20975 -9670
rect 12987 -10493 13203 -10489
rect 17884 -10525 20975 -10431
rect 17884 -10527 18819 -10525
rect 21051 -10626 21142 -9591
rect 21212 -10020 21271 -9333
rect 21443 -9335 21453 -9333
rect 21591 -9335 21601 -9042
rect 21447 -9347 21597 -9335
rect 20709 -10627 21142 -10626
rect 20709 -10737 21342 -10627
rect 20709 -10769 21343 -10737
rect 18208 -10967 18288 -10955
rect 18373 -10967 18743 -10965
rect 10106 -13570 17240 -11056
rect 18208 -11383 18214 -10967
rect 18282 -11383 18743 -10967
rect 18208 -11394 18743 -11383
rect 18208 -11395 18288 -11394
rect 18833 -11398 19211 -10955
rect 19303 -11398 19681 -10955
rect 19772 -11392 20150 -10949
rect 20236 -11398 20614 -10955
rect 20709 -11388 20852 -10769
rect 21142 -10966 21212 -10954
rect 21142 -10971 21148 -10966
rect 20949 -11371 21148 -10971
rect 21206 -11371 21212 -10966
rect 20949 -11383 21212 -11371
rect 20949 -11405 21206 -11383
rect 10106 -13678 13910 -13570
rect 10106 -13709 13209 -13678
rect 13259 -13709 13910 -13678
rect 10106 -13938 13910 -13709
rect 10106 -14138 12808 -13938
rect 13008 -14138 13910 -13938
rect 10106 -14386 13910 -14138
rect 14002 -13940 14626 -13659
rect 14002 -14142 14206 -13940
rect 14408 -14142 14626 -13940
rect 14002 -14303 14626 -14142
rect 14723 -14386 17240 -13570
rect 10106 -16903 17240 -14386
rect 18148 -11613 18331 -11597
rect 18148 -12031 18214 -11613
rect 18272 -12031 18514 -11613
rect 18148 -12050 18514 -12031
rect 18605 -12044 18983 -11601
rect 19074 -12050 19452 -11607
rect 19544 -12050 19922 -11607
rect 20007 -12050 20385 -11607
rect 20477 -12050 20855 -11607
rect 21154 -11611 21224 -11599
rect 21154 -11622 21160 -11611
rect 20943 -12016 21160 -11622
rect 21218 -12016 21224 -11611
rect 20943 -12022 21224 -12016
rect 21154 -12028 21224 -12022
rect 18148 -13676 18331 -12050
rect 21253 -12359 21343 -10769
rect 20940 -12449 21343 -12359
rect 19420 -12533 20075 -12527
rect 19420 -12679 19432 -12533
rect 20063 -12679 20075 -12533
rect 19420 -12685 20075 -12679
rect 19461 -12845 20035 -12685
rect 18680 -12858 20792 -12845
rect 18680 -12892 19251 -12858
rect 20235 -12892 20792 -12858
rect 18680 -12939 20792 -12892
rect 18680 -12951 20795 -12939
rect 18680 -13127 18697 -12951
rect 18731 -13127 20755 -12951
rect 20789 -13127 20795 -12951
rect 18680 -13139 20795 -13127
rect 18680 -13186 20792 -13139
rect 18680 -13220 19251 -13186
rect 20235 -13220 20792 -13186
rect 18680 -13222 20792 -13220
rect 19239 -13226 20247 -13222
rect 20940 -13364 21091 -12449
rect 19704 -13515 21091 -13364
rect 19704 -13601 19855 -13515
rect 21650 -13565 21815 -13559
rect 18148 -13695 18768 -13676
rect 18148 -15280 18779 -13695
rect 18148 -18059 18331 -15280
rect 18646 -15290 18779 -15280
rect 19279 -15337 20279 -13601
rect 20773 -13730 21650 -13565
rect 20773 -14079 20938 -13730
rect 21650 -13736 21815 -13730
rect 20773 -14091 20946 -14079
rect 20773 -14582 20883 -14091
rect 20940 -14582 20946 -14091
rect 20773 -14594 20946 -14582
rect 20773 -15297 20938 -14594
rect 18682 -16123 20794 -15746
rect 19439 -16295 20013 -16123
rect 19399 -16301 20054 -16295
rect 19399 -16447 19411 -16301
rect 20042 -16447 20054 -16301
rect 19399 -16453 20054 -16447
rect 18033 -18071 18391 -18059
rect 18033 -18727 18039 -18071
rect 18385 -18727 18391 -18071
rect 18033 -18739 18391 -18727
<< via1 >>
rect 12751 -5827 12822 -5607
rect 13085 -5829 13156 -5609
rect 13747 -5831 13818 -5611
rect 14080 -5832 14151 -5612
rect 14409 -5927 14481 -5618
rect 12751 -6648 12829 -6212
rect 13085 -6643 13156 -6423
rect 13419 -6644 13490 -6424
rect 14081 -6645 14152 -6425
rect 14413 -6645 14484 -6425
rect 9162 -7899 9256 -7804
rect 8056 -8200 8192 -7943
rect 10168 -8200 10304 -7941
rect 16342 -7318 16464 -7196
rect 9175 -8707 9245 -8453
rect 14500 -8272 14584 -8188
rect 16807 -7318 16929 -7196
rect 12783 -8562 12847 -8289
rect 17518 -8462 17574 -8335
rect 10708 -9018 10936 -8790
rect 12808 -9012 12968 -8816
rect 17365 -8788 17417 -8736
rect 14206 -9011 14407 -8810
rect 12808 -9017 12908 -9012
rect 14500 -9200 14584 -9116
rect 12238 -9657 12466 -9429
rect 12808 -9734 12908 -9634
rect 12811 -10469 12899 -10157
rect 18832 -8892 20522 -8838
rect 18096 -9331 18226 -9060
rect 13433 -10169 13608 -9994
rect 17135 -10169 17310 -9994
rect 19295 -9796 19405 -9650
rect 18909 -10169 19084 -9994
rect 20240 -9792 20359 -9659
rect 20494 -10169 20669 -9994
rect 21453 -9335 21591 -9042
rect 12808 -14138 13008 -13938
rect 14206 -14142 14408 -13940
rect 19432 -12679 20063 -12533
rect 21650 -13730 21815 -13565
rect 19411 -16447 20042 -16301
<< metal2 >>
rect 14412 -5365 15123 -5295
rect 12751 -5607 12822 -5597
rect 13085 -5607 13156 -5599
rect 12822 -5609 13156 -5607
rect 12822 -5827 13085 -5609
rect 12751 -5828 13085 -5827
rect 12751 -5837 12822 -5828
rect 13085 -5839 13156 -5829
rect 13747 -5611 13818 -5601
rect 14080 -5611 14151 -5602
rect 14412 -5608 14482 -5365
rect 13818 -5612 14151 -5611
rect 13818 -5831 14080 -5612
rect 13747 -5832 14080 -5831
rect 13747 -5841 13818 -5832
rect 14080 -5842 14151 -5832
rect 14409 -5618 14482 -5608
rect 14481 -5927 14482 -5618
rect 14409 -5937 14482 -5927
rect 14412 -6044 14482 -5937
rect 12751 -6212 12829 -6202
rect 12751 -6658 12829 -6648
rect 13085 -6421 13156 -6413
rect 13419 -6421 13490 -6414
rect 13085 -6423 13491 -6421
rect 14081 -6423 14152 -6415
rect 14413 -6423 14484 -6415
rect 13156 -6424 13491 -6423
rect 13156 -6642 13419 -6424
rect 13085 -6653 13156 -6643
rect 13490 -6642 13491 -6424
rect 14080 -6425 14484 -6423
rect 14080 -6644 14081 -6425
rect 13419 -6654 13490 -6644
rect 14152 -6644 14413 -6425
rect 14081 -6655 14152 -6645
rect 14413 -6655 14484 -6645
rect 12755 -6973 12824 -6658
rect 12755 -7042 12969 -6973
rect 15053 -6976 15123 -5365
rect 9162 -7804 9256 -7794
rect 9162 -7909 9256 -7899
rect 8056 -7943 8192 -7933
rect 8056 -8210 8192 -8200
rect 9169 -8283 9253 -7909
rect 10168 -7941 10304 -7931
rect 10168 -8210 10304 -8200
rect 12783 -8283 12847 -8279
rect 9169 -8289 12852 -8283
rect 9169 -8453 12783 -8289
rect 9169 -8707 9175 -8453
rect 9245 -8562 12783 -8453
rect 12847 -8562 12852 -8289
rect 9245 -8575 12852 -8562
rect 9245 -8707 9253 -8575
rect 9169 -8749 9253 -8707
rect 10702 -9018 10708 -8790
rect 10936 -9018 10942 -8790
rect 12900 -8810 12969 -7042
rect 14271 -7046 15123 -6976
rect 14271 -8804 14341 -7046
rect 16807 -7196 16929 -7190
rect 16336 -7318 16342 -7196
rect 16464 -7318 16807 -7196
rect 16807 -7324 16929 -7318
rect 14500 -8188 14584 -8182
rect 12808 -8816 12969 -8810
rect 12968 -8989 12969 -8816
rect 14206 -8810 14407 -8804
rect 12908 -9017 12968 -9012
rect 10708 -9429 10936 -9018
rect 12808 -9022 12968 -9017
rect 14500 -8830 14584 -8272
rect 17523 -8325 17566 -8323
rect 17518 -8335 17574 -8325
rect 17518 -8472 17574 -8462
rect 17359 -8788 17365 -8736
rect 17417 -8741 17423 -8736
rect 17523 -8741 17566 -8472
rect 17417 -8784 17566 -8741
rect 17417 -8788 17423 -8784
rect 17523 -8796 17566 -8784
rect 18832 -8830 20522 -8828
rect 14496 -8838 21815 -8830
rect 14496 -8892 18832 -8838
rect 20522 -8892 21815 -8838
rect 14496 -8995 21815 -8892
rect 12808 -9061 12908 -9022
rect 12797 -9236 13608 -9061
rect 14206 -9198 14407 -9011
rect 10708 -9657 12238 -9429
rect 12466 -9657 12472 -9429
rect 12808 -9634 12908 -9236
rect 12808 -9740 12908 -9734
rect 13433 -9994 13608 -9236
rect 14204 -9389 14407 -9198
rect 14500 -9116 14584 -8995
rect 21453 -9042 21591 -9032
rect 14500 -9206 14584 -9200
rect 18096 -9060 18226 -9050
rect 18096 -9341 18226 -9331
rect 21453 -9345 21591 -9335
rect 14204 -9574 20367 -9389
rect 14204 -9607 20372 -9574
rect 12811 -10157 12899 -10147
rect 13433 -10175 13608 -10169
rect 12811 -10479 12899 -10469
rect 12819 -10762 12891 -10479
rect 14206 -10749 14407 -9607
rect 14495 -9613 20372 -9607
rect 19286 -9650 19423 -9613
rect 19286 -9685 19295 -9650
rect 19405 -9685 19423 -9650
rect 20235 -9659 20372 -9613
rect 19295 -9806 19405 -9796
rect 20240 -9802 20359 -9792
rect 17135 -9994 17310 -9988
rect 17310 -10169 18909 -9994
rect 19084 -10169 20494 -9994
rect 20669 -10169 20675 -9994
rect 17135 -10175 17310 -10169
rect 12808 -10930 13009 -10762
rect 12808 -13938 13008 -10930
rect 12808 -14144 13008 -14138
rect 14206 -13940 14408 -10749
rect 19432 -12533 20063 -12523
rect 19432 -12689 20063 -12679
rect 21650 -13565 21815 -8995
rect 21644 -13730 21650 -13565
rect 21815 -13730 21821 -13565
rect 14206 -14148 14408 -14142
rect 19411 -16301 20042 -16291
rect 19411 -16457 20042 -16447
<< via2 >>
rect 8056 -8200 8192 -7943
rect 10168 -8200 10304 -7941
rect 18096 -9331 18226 -9060
rect 21453 -9335 21591 -9042
rect 19432 -12679 20063 -12533
rect 19411 -16447 20042 -16301
<< metal3 >>
rect 8010 -5154 18268 -4940
rect 8010 -7943 8224 -5154
rect 8010 -8200 8056 -7943
rect 8192 -8200 8224 -7943
rect 8010 -8214 8224 -8200
rect 10114 -7941 10328 -5154
rect 10114 -8200 10168 -7941
rect 10304 -8200 10328 -7941
rect 10114 -8290 10328 -8200
rect 18054 -7660 18268 -5154
rect 18054 -7874 21624 -7660
rect 18054 -9060 18268 -7874
rect 18054 -9331 18096 -9060
rect 18226 -9331 18268 -9060
rect 18054 -12483 18268 -9331
rect 21410 -9042 21624 -7874
rect 21410 -9335 21453 -9042
rect 21591 -9335 21624 -9042
rect 21410 -9448 21624 -9335
rect 18054 -12533 20125 -12483
rect 18054 -12679 19432 -12533
rect 20063 -12679 20125 -12533
rect 18054 -12697 20125 -12679
rect 18073 -16274 18287 -12697
rect 18073 -16301 20075 -16274
rect 18073 -16447 19411 -16301
rect 20042 -16447 20075 -16301
rect 18073 -16488 20075 -16447
use sky130_fd_pr__nfet_01v8_lvt_63HJ42  sky130_fd_pr__nfet_01v8_lvt_63HJ42_0
timestamp 1724943425
transform 1 0 17310 0 1 -8541
box -424 -257 424 257
use sky130_fd_pr__nfet_01v8_lvt_JQYUHL  sky130_fd_pr__nfet_01v8_lvt_JQYUHL_0
timestamp 1725314430
transform 1 0 13682 0 1 -7939
box -2603 -857 2603 857
use sky130_fd_pr__pfet_01v8_lvt_9BX3CZ  sky130_fd_pr__pfet_01v8_lvt_9BX3CZ_0
timestamp 1725314430
transform 1 0 9212 0 1 -8289
box -839 -498 839 464
use sky130_fd_pr__pfet_01v8_lvt_66XZ34  sky130_fd_pr__pfet_01v8_lvt_66XZ34_0
timestamp 1725402679
transform 1 0 19817 0 1 -9477
box -1487 -598 1487 564
use sky130_fd_pr__pfet_01v8_lvt_AZ5TEV  sky130_fd_pr__pfet_01v8_lvt_AZ5TEV_0
timestamp 1725483475
transform 1 0 19731 0 1 -15929
box -1094 -200 1094 200
use sky130_fd_pr__pfet_01v8_lvt_AZ5TEV  sky130_fd_pr__pfet_01v8_lvt_AZ5TEV_1
timestamp 1725483475
transform -1 0 19743 0 -1 -13039
box -1094 -200 1094 200
use sky130_fd_pr__pfet_01v8_lvt_W4537V  sky130_fd_pr__pfet_01v8_lvt_W4537V_0
timestamp 1725483475
transform 1 0 19778 0 1 -14479
box -1196 -973 1196 973
use sky130_fd_pr__res_xhigh_po_0p35_9LVS8Q  sky130_fd_pr__res_xhigh_po_0p35_9LVS8Q_0
timestamp 1725526980
transform -1 0 14281 0 -1 -6128
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p35_32GTF4  sky130_fd_pr__res_xhigh_po_0p35_32GTF4_0
timestamp 1725527848
transform -1 0 12858 0 -1 -9950
box -367 -687 367 687
use sky130_fd_pr__res_xhigh_po_0p35_ZJVS8Y  sky130_fd_pr__res_xhigh_po_0p35_ZJVS8Y_0
timestamp 1725526980
transform -1 0 12956 0 -1 -6128
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p69_5SXZXT  sky130_fd_pr__res_xhigh_po_0p69_5SXZXT_0
timestamp 1725054543
transform 1 0 19728 0 1 -11508
box -1522 -708 1522 708
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2 ~/pdk/sky130A/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 5 1288
timestamp 1704896540
transform 0 -1 17563 1 0 -17226
box 0 0 1340 1340
<< labels >>
rlabel metal2 17523 -8789 17566 -8724 1 Gcm2
rlabel metal2 9266 -8510 9385 -8302 1 Gcm1
rlabel metal1 17170 -7775 17273 -7598 1 Sop
flabel metal3 10099 -5094 10407 -4946 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel psubdiffcont 23115 -4597 23922 -3277 0 FreeSans 160 0 0 0 VSS
port 3 nsew
rlabel metal1 12209 -8994 12528 -8798 1 PLUS
rlabel metal1 13844 -8986 14131 -8814 1 MINUS
flabel metal1 20919 -10749 21242 -10637 0 FreeSans 160 0 0 0 Vbgr
port 2 nsew
flabel metal1 10696 -6750 10856 -6430 0 FreeSans 160 0 0 0 VSS
port 3 nsew
<< end >>
