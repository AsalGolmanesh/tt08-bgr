* NGSPICE file created from core_prel_parax.ext - technology: sky130A

.subckt core_prel_parax VDD Vbgr VSS
X0 VDD.t17 w_21453_n6696.t13 a_17750_n8805.t2 VDD.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 Gcm2 w_21453_n6696.t14 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_17750_n8805.t3 XQ2[0|0].Emitter VSS.t79 sky130_fd_pr__res_xhigh_po_0p35 l=0.9
X3 VSS.t78 VSS.t75 VSS.t77 VSS.t76 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X4 VSS.t1 a_23542_n10376# VSS.t0 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X5 VDD.t32 VDD.t30 w_21453_n6696.t0 VDD.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X6 MINUS.t2 w_21453_n6696.t15 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X7 VSS.t38 VSS.t74 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X8 VSS.t40 VSS.t73 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X9 VSS.t44 VSS.t72 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X10 w_21453_n6696.t5 VDD.t27 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X11 w_21453_n6696.t3 a_17692_n8717.t8 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X12 a_25081_n8277# a_25579_n8877# VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X13 Vbgr.t0 a_25414_n10376# VSS.t6 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X14 VSS.t38 VSS.t71 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X15 VSS.t40 VSS.t70 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X16 VSS.t40 VSS.t69 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X17 VDD.t11 w_21453_n6696.t16 Vbgr.t2 VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X18 VSS.t68 VSS.t66 a_17692_n8717.t1 VSS.t67 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=4
X19 VSS.t17 VSS.t18 VSS.t16 sky130_fd_pr__res_xhigh_po_0p35 l=1
X20 Gcm2 Gcm2 VSS.t25 VSS.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X21 VSS.t38 VSS.t60 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X22 VSS.t42 VSS.t65 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X23 VSS.t64 VSS.t62 Gcm2 VSS.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X24 VSS.t31 VSS.t59 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X25 VSS.t31 VSS.t58 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X26 VSS.t31 VSS.t61 MINUS.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X27 a_25180_n9724# a_25414_n10376# VSS.t6 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X28 VSS.t15 a_23825_n8877# VSS.t14 sky130_fd_pr__res_xhigh_po_0p35 l=1
X29 VSS.t33 VSS.t57 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X30 VSS.t42 VSS.t56 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X31 a_24157_n8277# a_24323_n8877# VSS.t13 sky130_fd_pr__res_xhigh_po_0p35 l=1
X32 VSS.t4 VSS.t5 VSS.t3 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X33 VDD.t26 VDD.t24 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=0.5
X34 a_23991_n8277# a_24915_n8877# VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X35 VSS.t44 VSS.t55 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X36 VSS.t42 VSS.t54 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X37 VSS.t42 VSS.t53 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X38 VDD.t9 w_21453_n6696.t17 Gcm2 VDD.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X39 VDD.t7 w_21453_n6696.t18 MINUS.t1 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X40 w_21453_n6696.t4 MINUS.t4 Sop.t5 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X41 a_25247_n8277# MINUS.t0 VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X42 a_24712_n9724# a_24946_n10376# VSS.t6 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X43 VSS.t33 VSS.t52 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X44 VSS.t33 VSS.t51 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X45 VSS.t33 VSS.t50 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X46 w_21453_n6696.t7 Vbgr.t3 VSS.t80 w_21453_n6696.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X47 a_23493_n8277# VSS.t88 VSS.t87 sky130_fd_pr__res_xhigh_po_0p35 l=1
X48 a_23493_n8277# a_23659_n8877# VSS.t11 sky130_fd_pr__res_xhigh_po_0p35 l=1
X49 VSS.t40 VSS.t49 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X50 VSS.t44 VSS.t48 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X51 w_21453_n6696.t2 Vbgr.t4 VSS.t19 w_21453_n6696.t1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X52 Sop.t3 a_17750_n8805.t4 a_17692_n8717.t6 VSS.t83 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X53 a_24157_n8277# a_23659_n8877# VSS.t89 sky130_fd_pr__res_xhigh_po_0p35 l=1
X54 VSS.t9 VSS.t10 VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X55 a_24244_n9724# a_24478_n10376# VSS.t7 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X56 a_24712_n9724# a_24478_n10376# VSS.t6 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X57 VSS.t38 VSS.t47 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X58 w_21453_n6696.t10 Vbgr.t5 VSS.t84 w_21453_n6696.t9 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X59 a_17750_n8805.t1 w_21453_n6696.t19 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X60 VSS.t31 VSS.t46 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X61 VDD.t36 a_17692_n8717.t9 w_21453_n6696.t8 VDD.t35 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X62 VDD.t23 VDD.t20 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.5
X63 a_23991_n8277# a_23825_n8877# VSS.t28 sky130_fd_pr__res_xhigh_po_0p35 l=1
X64 a_25081_n8277# a_24915_n8877# VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X65 a_25247_n8277# a_24323_n8877# VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X66 Sop.t1 Gcm2 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X67 a_24244_n9724# a_24010_n10376# VSS.t2 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X68 VSS.t44 VSS.t45 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X69 VSS.t44 VSS.t43 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X70 w_21453_n6696.t12 Vbgr.t6 VSS.t86 w_21453_n6696.t11 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X71 VSS.t21 Gcm2 Sop.t0 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X72 Sop.t4 MINUS.t5 w_21453_n6696.t4 VSS.t85 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X73 VSS.t26 VSS.t27 VSS.t6 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X74 a_23776_n9724# a_24010_n10376# VSS.t12 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X75 VSS.t42 VSS.t41 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X76 VDD.t34 a_17692_n8717.t4 a_17692_n8717.t5 VDD.t33 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X77 a_17692_n8717.t7 a_17750_n8805.t5 Sop.t2 VSS.t82 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X78 a_17750_n8805.t0 a_25579_n8877# VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1
X79 a_17692_n8717.t3 a_17692_n8717.t2 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X80 Vbgr.t1 w_21453_n6696.t20 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X81 VSS.t40 VSS.t39 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X82 VSS.t38 VSS.t37 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X83 a_17692_n8717.t0 VSS.t34 VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=4
X84 a_23776_n9724# a_23542_n10376# VSS.t81 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X85 VSS.t33 VSS.t32 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X86 VSS.t31 VSS.t30 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X87 a_25180_n9724# a_24946_n10376# VSS.t6 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
R0 w_21453_n6696.n0 w_21453_n6696.t16 674.212
R1 w_21453_n6696.n0 w_21453_n6696.t14 674.149
R2 w_21453_n6696.n0 w_21453_n6696.t17 674.149
R3 w_21453_n6696.n0 w_21453_n6696.t19 674.149
R4 w_21453_n6696.n0 w_21453_n6696.t13 674.149
R5 w_21453_n6696.n0 w_21453_n6696.t15 674.149
R6 w_21453_n6696.n0 w_21453_n6696.t18 674.149
R7 w_21453_n6696.n0 w_21453_n6696.t20 674.149
R8 w_21453_n6696.n0 w_21453_n6696.t2 228.215
R9 w_21453_n6696.n0 w_21453_n6696.t7 228.215
R10 w_21453_n6696.n0 w_21453_n6696.t12 228.215
R11 w_21453_n6696.n0 w_21453_n6696.t10 228.215
R12 w_21453_n6696.n1 w_21453_n6696.t4 210.763
R13 w_21453_n6696.t6 w_21453_n6696.t1 173.161
R14 w_21453_n6696.t11 w_21453_n6696.t9 173.161
R15 w_21453_n6696.n1 w_21453_n6696.n2 153.768
R16 w_21453_n6696.n4 w_21453_n6696.n1 152.613
R17 w_21453_n6696.n3 w_21453_n6696.t6 86.5808
R18 w_21453_n6696.n3 w_21453_n6696.t11 86.5808
R19 w_21453_n6696.n0 w_21453_n6696.n3 17.8715
R20 w_21453_n6696.n1 w_21453_n6696.n0 9.42554
R21 w_21453_n6696.n2 w_21453_n6696.t8 7.14175
R22 w_21453_n6696.n2 w_21453_n6696.t5 7.14175
R23 w_21453_n6696.t0 w_21453_n6696.n4 7.14175
R24 w_21453_n6696.n4 w_21453_n6696.t3 7.14175
R25 a_17750_n8805.n2 a_17750_n8805.n0 276.264
R26 a_17750_n8805.n1 a_17750_n8805.t4 68.6435
R27 a_17750_n8805.n1 a_17750_n8805.t5 66.1962
R28 a_17750_n8805.n3 a_17750_n8805.t3 53.4029
R29 a_17750_n8805.t0 a_17750_n8805.n3 43.7745
R30 a_17750_n8805.n2 a_17750_n8805.n1 16.4639
R31 a_17750_n8805.n0 a_17750_n8805.t2 2.857
R32 a_17750_n8805.n0 a_17750_n8805.t1 2.857
R33 a_17750_n8805.n3 a_17750_n8805.n2 0.394995
R34 VDD.n11 VDD.t24 675.381
R35 VDD.n22 VDD.t20 674.89
R36 VDD.n24 VDD.t23 278.337
R37 VDD.t26 VDD.n10 278.334
R38 VDD.n21 VDD.n20 275.077
R39 VDD.n19 VDD.n18 275.077
R40 VDD.n17 VDD.n16 275.077
R41 VDD.n15 VDD.n14 275.077
R42 VDD.n13 VDD.n12 275.077
R43 VDD.t28 VDD.n33 271.897
R44 VDD.n8 VDD.t31 257.913
R45 VDD.n6 VDD.t30 192.475
R46 VDD.n1 VDD.t27 192.475
R47 VDD.n27 VDD.n26 162.465
R48 VDD.n7 VDD.t32 159.048
R49 VDD.n0 VDD.t29 159.048
R50 VDD.t31 VDD.t18 152.52
R51 VDD.t18 VDD.t33 152.52
R52 VDD.t0 VDD.t35 152.52
R53 VDD.t35 VDD.t28 152.52
R54 VDD.n25 VDD.n23 152.345
R55 VDD.n3 VDD.n2 151.905
R56 VDD.n5 VDD.n4 151.905
R57 VDD.t21 VDD.n25 143.857
R58 VDD.n26 VDD.t25 140.78
R59 VDD.n26 VDD.n10 118.692
R60 VDD.n25 VDD.n24 116.584
R61 VDD VDD.t33 98.1337
R62 VDD.t25 VDD.t10 69.427
R63 VDD.t10 VDD.t2 69.427
R64 VDD.t2 VDD.t6 69.427
R65 VDD.t6 VDD.t12 69.427
R66 VDD.t12 VDD.t16 69.427
R67 VDD.t16 VDD.t4 69.427
R68 VDD.t4 VDD.t8 69.427
R69 VDD.t8 VDD.t14 69.427
R70 VDD.t14 VDD.t21 69.427
R71 VDD VDD.t0 54.3876
R72 VDD.n2 VDD.t1 7.14175
R73 VDD.n2 VDD.t36 7.14175
R74 VDD.n4 VDD.t19 7.14175
R75 VDD.n4 VDD.t34 7.14175
R76 VDD.n20 VDD.t15 2.857
R77 VDD.n20 VDD.t22 2.857
R78 VDD.n18 VDD.t5 2.857
R79 VDD.n18 VDD.t9 2.857
R80 VDD.n16 VDD.t13 2.857
R81 VDD.n16 VDD.t17 2.857
R82 VDD.n14 VDD.t3 2.857
R83 VDD.n14 VDD.t7 2.857
R84 VDD.n12 VDD.t26 2.857
R85 VDD.n12 VDD.t11 2.857
R86 VDD.n23 VDD.n9 2.26217
R87 VDD.n28 VDD.n27 2.26217
R88 VDD.n33 VDD.n32 2.20468
R89 VDD.n28 VDD.n10 2.09911
R90 VDD.n24 VDD.n9 1.99684
R91 VDD.n32 VDD.n8 1.2782
R92 VDD.n30 VDD.n29 0.975785
R93 VDD.n29 VDD.n28 0.723704
R94 VDD.n5 VDD.n3 0.233352
R95 VDD.n29 VDD.n9 0.218658
R96 VDD.n3 VDD.n1 0.164385
R97 VDD.n6 VDD.n5 0.164385
R98 VDD.n22 VDD.n21 0.143692
R99 VDD.n13 VDD.n11 0.1405
R100 VDD.n15 VDD.n13 0.122038
R101 VDD.n17 VDD.n15 0.122038
R102 VDD.n19 VDD.n17 0.122038
R103 VDD.n21 VDD.n19 0.122038
R104 VDD.n33 VDD.n0 0.0940792
R105 VDD.n8 VDD.n7 0.086224
R106 VDD.n1 VDD.n0 0.0445574
R107 VDD.n7 VDD.n6 0.0445574
R108 VDD.n30 VDD 0.0299078
R109 VDD VDD.n31 0.024
R110 VDD.n31 VDD 0.023873
R111 VDD.n32 VDD 0.0176141
R112 VDD.n31 VDD.n30 0.00558108
R113 VDD.n23 VDD.n22 0.00176918
R114 VDD.n27 VDD.n11 0.00165385
R115 VSS.n1874 VSS.n1870 20051.4
R116 VSS.n1891 VSS.n1870 16174.6
R117 VSS.n4639 VSS.n1393 12208.2
R118 VSS.n1899 VSS.n1870 9706.76
R119 VSS.n4625 VSS.n1402 7289
R120 VSS.n4626 VSS.n1402 7289
R121 VSS.n4663 VSS.n1369 7289
R122 VSS.n4658 VSS.n1369 7289
R123 VSS.n1378 VSS.n1370 6993.5
R124 VSS.n4620 VSS.n1401 6993.5
R125 VSS.n4153 VSS.n1899 4974.74
R126 VSS.n4626 VSS.n1401 3743
R127 VSS.n4658 VSS.n1378 3743
R128 VSS.n4625 VSS.n4620 3644.5
R129 VSS.n4663 VSS.n1370 3644.5
R130 VSS.n4154 VSS.n4153 3409.8
R131 VSS.n4155 VSS.t38 2890.74
R132 VSS.n4182 VSS.n4180 2277.04
R133 VSS.n4072 VSS.n4071 1851.56
R134 VSS.n4729 VSS.n4728 1851.56
R135 VSS.n4708 VSS.n4707 1851.56
R136 VSS.n1684 VSS.n1683 1801.72
R137 VSS.n4986 VSS.n4985 1801.72
R138 VSS.n675 VSS.n674 1801.72
R139 VSS.n2625 VSS.n2589 1634.59
R140 VSS.n2789 VSS.n2788 1559.06
R141 VSS.n2788 VSS.n2787 1559.06
R142 VSS.n2787 VSS.n2761 1559.06
R143 VSS.n2781 VSS.n2761 1559.06
R144 VSS.n2781 VSS.n2780 1559.06
R145 VSS.n2777 VSS.n2776 1559.06
R146 VSS.n2776 VSS.n2775 1559.06
R147 VSS.n2775 VSS.n2766 1559.06
R148 VSS.n2768 VSS.n2766 1559.06
R149 VSS.n2768 VSS.n2767 1559.06
R150 VSS.n4071 VSS.n4070 1559.06
R151 VSS.n4070 VSS.n4001 1559.06
R152 VSS.n4064 VSS.n4001 1559.06
R153 VSS.n4064 VSS.n1172 1559.06
R154 VSS.n4007 VSS.n1173 1559.06
R155 VSS.n4057 VSS.n4007 1559.06
R156 VSS.n4057 VSS.n4056 1559.06
R157 VSS.n4056 VSS.n4055 1559.06
R158 VSS.n4055 VSS.n1174 1559.06
R159 VSS.n4728 VSS.n4727 1559.06
R160 VSS.n4727 VSS.n1167 1559.06
R161 VSS.n1171 VSS.n1167 1559.06
R162 VSS.n4720 VSS.n1171 1559.06
R163 VSS.n3907 VSS.n1175 1559.06
R164 VSS.n3913 VSS.n3907 1559.06
R165 VSS.n3914 VSS.n3913 1559.06
R166 VSS.n3915 VSS.n3914 1559.06
R167 VSS.n3915 VSS.n1176 1559.06
R168 VSS.n1683 VSS.n1655 1559.06
R169 VSS.n1677 VSS.n1655 1559.06
R170 VSS.n1677 VSS.n1676 1559.06
R171 VSS.n1673 VSS.n1672 1559.06
R172 VSS.n1672 VSS.n1671 1559.06
R173 VSS.n1671 VSS.n1660 1559.06
R174 VSS.n1665 VSS.n1660 1559.06
R175 VSS.n1665 VSS.n1664 1559.06
R176 VSS.n4985 VSS.n766 1559.06
R177 VSS.n4979 VSS.n766 1559.06
R178 VSS.n4979 VSS.n4978 1559.06
R179 VSS.n4975 VSS.n4974 1559.06
R180 VSS.n4974 VSS.n4973 1559.06
R181 VSS.n4973 VSS.n771 1559.06
R182 VSS.n4967 VSS.n771 1559.06
R183 VSS.n4967 VSS.n4966 1559.06
R184 VSS.n674 VSS.n646 1559.06
R185 VSS.n668 VSS.n646 1559.06
R186 VSS.n668 VSS.n667 1559.06
R187 VSS.n664 VSS.n663 1559.06
R188 VSS.n663 VSS.n662 1559.06
R189 VSS.n662 VSS.n651 1559.06
R190 VSS.n656 VSS.n651 1559.06
R191 VSS.n656 VSS.n655 1559.06
R192 VSS.n4707 VSS.n4706 1559.06
R193 VSS.n4706 VSS.n1210 1559.06
R194 VSS.n1211 VSS.n1210 1559.06
R195 VSS.n1211 VSS.n1177 1559.06
R196 VSS.n4697 VSS.n1178 1559.06
R197 VSS.n4697 VSS.n4696 1559.06
R198 VSS.n4696 VSS.n4695 1559.06
R199 VSS.n4695 VSS.n1216 1559.06
R200 VSS.n1216 VSS.n1179 1559.06
R201 VSS.n4163 VSS.n1866 1540.86
R202 VSS.n4164 VSS.n4163 1540.86
R203 VSS.n4165 VSS.n4164 1540.86
R204 VSS.n4172 VSS.n1862 1540.86
R205 VSS.n4173 VSS.n4172 1540.86
R206 VSS.n4174 VSS.n4173 1540.86
R207 VSS.n4174 VSS.n1859 1540.86
R208 VSS.n4178 VSS.n1859 1540.86
R209 VSS.n4179 VSS.n4178 1540.86
R210 VSS.n4183 VSS.n4182 1540.86
R211 VSS.n4208 VSS.n4183 1540.86
R212 VSS.n4208 VSS.n4207 1540.86
R213 VSS.n4207 VSS.n4206 1540.86
R214 VSS.n4206 VSS.n1183 1540.86
R215 VSS.n4199 VSS.n1184 1540.86
R216 VSS.n4199 VSS.n4198 1540.86
R217 VSS.n4198 VSS.n4197 1540.86
R218 VSS.n4197 VSS.n4187 1540.86
R219 VSS.n4191 VSS.n4187 1540.86
R220 VSS.n5370 VSS.n165 1497.55
R221 VSS.n4637 VSS.n4634 1332.39
R222 VSS.n1397 VSS.n1394 1311.29
R223 VSS.n4180 VSS.n4179 1284.05
R224 VSS.t33 VSS.n1185 1103.21
R225 VSS.n2780 VSS.t38 1056.69
R226 VSS.t33 VSS.n1172 1056.69
R227 VSS.n4720 VSS.t33 1056.69
R228 VSS.n1676 VSS.t44 1056.69
R229 VSS.n4978 VSS.t44 1056.69
R230 VSS.n667 VSS.t44 1056.69
R231 VSS.t33 VSS.n1177 1056.69
R232 VSS.n4165 VSS.t38 1044.36
R233 VSS.t33 VSS.n1183 1044.36
R234 VSS.n5564 VSS.n5563 888.997
R235 VSS.n4618 VSS.n1378 857.529
R236 VSS.n4618 VSS.n1401 857.529
R237 VSS.n4180 VSS.n1857 855.557
R238 VSS.n2569 VSS.n1265 855.557
R239 VSS.n2545 VSS.n2389 855.557
R240 VSS.n4641 VSS.n1390 855.557
R241 VSS.n2286 VSS.n20 855.557
R242 VSS.n4619 VSS.n1370 840.148
R243 VSS.n4620 VSS.n4619 840.148
R244 VSS.n1898 VSS.n1897 829.587
R245 VSS.n1898 VSS.n1 827.635
R246 VSS.n5565 VSS.n5564 770.559
R247 VSS.n5566 VSS.n1 760.035
R248 VSS.n4153 VSS.n4152 728.679
R249 VSS.n1871 VSS.n2 723.712
R250 VSS.n4156 VSS.n4154 718.693
R251 VSS.n2756 VSS.n2034 665.731
R252 VSS.n3062 VSS.t38 665.731
R253 VSS.n3148 VSS.t38 665.731
R254 VSS.n3222 VSS.t38 665.731
R255 VSS.n2767 VSS.t38 658.269
R256 VSS.t33 VSS.n1174 658.269
R257 VSS.t33 VSS.n1176 658.269
R258 VSS.n1664 VSS.t44 658.269
R259 VSS.n4966 VSS.t44 658.269
R260 VSS.n655 VSS.t44 658.269
R261 VSS.t33 VSS.n1179 658.269
R262 VSS.n2794 VSS.n2034 648.096
R263 VSS.n3114 VSS.t38 648.096
R264 VSS.n3186 VSS.t38 648.096
R265 VSS.n4078 VSS.t38 648.096
R266 VSS.n2357 VSS.n2322 641.164
R267 VSS.t35 VSS.t83 627.736
R268 VSS.n4191 VSS.n1185 616.342
R269 VSS.t82 VSS.t67 611.785
R270 VSS.n5224 VSS.n334 585
R271 VSS.n5224 VSS.n5223 585
R272 VSS.n358 VSS.n342 585
R273 VSS.n5218 VSS.n358 585
R274 VSS.n5216 VSS.n5215 585
R275 VSS.n4963 VSS.n4962 585
R276 VSS.n4403 VSS.n326 585
R277 VSS.n5234 VSS.n326 585
R278 VSS.n4403 VSS.n327 585
R279 VSS.n5234 VSS.n327 585
R280 VSS.n4992 VSS.n325 585
R281 VSS.n5234 VSS.n325 585
R282 VSS.n4992 VSS.n328 585
R283 VSS.n5234 VSS.n328 585
R284 VSS.n5232 VSS.n324 585
R285 VSS.n5234 VSS.n324 585
R286 VSS.n5233 VSS.n5232 585
R287 VSS.n5234 VSS.n5233 585
R288 VSS.n2363 VSS.n209 585
R289 VSS.n5231 VSS.n329 585
R290 VSS.n5231 VSS.n5230 585
R291 VSS.n4991 VSS.n760 585
R292 VSS.n4991 VSS.n4990 585
R293 VSS.n4402 VSS.n1584 585
R294 VSS.n4402 VSS.n4401 585
R295 VSS.n4401 VSS.n209 585
R296 VSS.n4401 VSS.n1687 585
R297 VSS.n1687 VSS.n1584 585
R298 VSS.n1584 VSS.n211 585
R299 VSS.n4990 VSS.n4989 585
R300 VSS.n4990 VSS.n211 585
R301 VSS.n4989 VSS.n760 585
R302 VSS.n760 VSS.n211 585
R303 VSS.n5230 VSS.n5229 585
R304 VSS.n5230 VSS.n211 585
R305 VSS.n5229 VSS.n329 585
R306 VSS.n329 VSS.n211 585
R307 VSS.n5437 VSS.n74 585
R308 VSS.n5437 VSS.n5436 585
R309 VSS.n74 VSS.n72 585
R310 VSS.n5436 VSS.n72 585
R311 VSS.n3476 VSS.n77 585
R312 VSS.n5436 VSS.n77 585
R313 VSS.n3476 VSS.n78 585
R314 VSS.n5436 VSS.n78 585
R315 VSS.n359 VSS.n76 585
R316 VSS.n5436 VSS.n76 585
R317 VSS.n359 VSS.n79 585
R318 VSS.n5436 VSS.n79 585
R319 VSS.n2284 VSS.n23 585
R320 VSS.n965 VSS.n846 585
R321 VSS.n967 VSS.n846 585
R322 VSS.n3681 VSS.n3477 585
R323 VSS.n3679 VSS.n3477 585
R324 VSS.n3540 VSS.n1451 585
R325 VSS.n1451 VSS.n73 585
R326 VSS.n73 VSS.n23 585
R327 VSS.n73 VSS.n70 585
R328 VSS.n3540 VSS.n70 585
R329 VSS.n3540 VSS.n25 585
R330 VSS.n3680 VSS.n3679 585
R331 VSS.n3679 VSS.n25 585
R332 VSS.n3681 VSS.n3680 585
R333 VSS.n3681 VSS.n25 585
R334 VSS.n967 VSS.n966 585
R335 VSS.n967 VSS.n25 585
R336 VSS.n966 VSS.n965 585
R337 VSS.n965 VSS.n25 585
R338 VSS.n5434 VSS.n75 585
R339 VSS.n5436 VSS.n75 585
R340 VSS.n5435 VSS.n5434 585
R341 VSS.n5436 VSS.n5435 585
R342 VSS.n5433 VSS.n80 585
R343 VSS.n80 VSS.n23 585
R344 VSS.n5433 VSS.n5432 585
R345 VSS.n5432 VSS.n5431 585
R346 VSS.n5432 VSS.n25 585
R347 VSS.n5431 VSS.n80 585
R348 VSS.n5429 VSS.n5428 585
R349 VSS.n5236 VSS.n320 585
R350 VSS.n5234 VSS.n320 585
R351 VSS.n5236 VSS.n5235 585
R352 VSS.n5235 VSS.n5234 585
R353 VSS.n322 VSS.n321 585
R354 VSS.n322 VSS.n209 585
R355 VSS.n643 VSS.n321 585
R356 VSS.n678 VSS.n643 585
R357 VSS.n643 VSS.n211 585
R358 VSS.n678 VSS.n322 585
R359 VSS.n5251 VSS.n303 585
R360 VSS.n5007 VSS.n743 585
R361 VSS.n4418 VSS.n1567 585
R362 VSS.n1227 VSS.n1220 585
R363 VSS.n4719 VSS.n1192 585
R364 VSS.n1338 VSS.n1306 585
R365 VSS.n5044 VSS.n5014 585
R366 VSS.n4048 VSS.n4047 585
R367 VSS.n3903 VSS.n3870 585
R368 VSS.n4051 VSS.n4009 585
R369 VSS.n4009 VSS.n1182 585
R370 VSS.n4051 VSS.n4050 585
R371 VSS.n4050 VSS.n1182 585
R372 VSS.n3920 VSS.n3919 585
R373 VSS.n3919 VSS.n1182 585
R374 VSS.n3921 VSS.n3920 585
R375 VSS.n3921 VSS.n1182 585
R376 VSS.n1304 VSS.n1303 585
R377 VSS.n1304 VSS.n1182 585
R378 VSS.n1303 VSS.n1276 585
R379 VSS.n1276 VSS.n1182 585
R380 VSS.n4688 VSS.n1219 585
R381 VSS.n4688 VSS.n1182 585
R382 VSS.n1221 VSS.n1219 585
R383 VSS.n1221 VSS.n1182 585
R384 VSS.n2708 VSS.n2239 585
R385 VSS.n4685 VSS.n1223 585
R386 VSS.n4687 VSS.n1223 585
R387 VSS.n1341 VSS.n1275 585
R388 VSS.n1277 VSS.n1275 585
R389 VSS.n3922 VSS.n3867 585
R390 VSS.n3868 VSS.n3867 585
R391 VSS.n4011 VSS.n4010 585
R392 VSS.n4013 VSS.n4010 585
R393 VSS.n4681 VSS.n1357 585
R394 VSS.n4681 VSS.n4680 585
R395 VSS.n4681 VSS.n1060 585
R396 VSS.n4014 VSS.n4013 585
R397 VSS.n4013 VSS.n1060 585
R398 VSS.n4014 VSS.n4011 585
R399 VSS.n4011 VSS.n1060 585
R400 VSS.n3923 VSS.n3868 585
R401 VSS.n3868 VSS.n1060 585
R402 VSS.n3923 VSS.n3922 585
R403 VSS.n3922 VSS.n1060 585
R404 VSS.n1340 VSS.n1277 585
R405 VSS.n1277 VSS.n1060 585
R406 VSS.n1341 VSS.n1340 585
R407 VSS.n1341 VSS.n1060 585
R408 VSS.n4687 VSS.n4686 585
R409 VSS.n4687 VSS.n1060 585
R410 VSS.n4686 VSS.n4685 585
R411 VSS.n4685 VSS.n1060 585
R412 VSS.n2709 VSS.n2708 585
R413 VSS.n2708 VSS.n1060 585
R414 VSS.n2791 VSS.n2037 585
R415 VSS.n2791 VSS.n2790 585
R416 VSS.n3065 VSS.n1994 585
R417 VSS.n3098 VSS.n1994 585
R418 VSS.n3097 VSS.n3065 585
R419 VSS.n3098 VSS.n3097 585
R420 VSS.n3097 VSS.n3096 585
R421 VSS.n3151 VSS.n1960 585
R422 VSS.n3183 VSS.n1960 585
R423 VSS.n3182 VSS.n3151 585
R424 VSS.n3183 VSS.n3182 585
R425 VSS.n3182 VSS.n3181 585
R426 VSS.n1915 VSS.n1913 585
R427 VSS.n1915 VSS.n1911 585
R428 VSS.n4076 VSS.n1913 585
R429 VSS.n4076 VSS.n1911 585
R430 VSS.n4076 VSS.n4075 585
R431 VSS.n4711 VSS.n1205 585
R432 VSS.n4709 VSS.n1205 585
R433 VSS.n4715 VSS.n1195 585
R434 VSS.n1195 VSS.n1129 585
R435 VSS.n3096 VSS.n1195 585
R436 VSS.n4732 VSS.n1160 585
R437 VSS.n4730 VSS.n1160 585
R438 VSS.n3181 VSS.n1160 585
R439 VSS.n4074 VSS.n3972 585
R440 VSS.n4074 VSS.n4073 585
R441 VSS.n4075 VSS.n4074 585
R442 VSS.n4073 VSS.n1199 585
R443 VSS.n4713 VSS.n1199 585
R444 VSS.n3972 VSS.n1200 585
R445 VSS.n4713 VSS.n1200 585
R446 VSS.n4730 VSS.n1165 585
R447 VSS.n4713 VSS.n1165 585
R448 VSS.n4732 VSS.n1158 585
R449 VSS.n4713 VSS.n1158 585
R450 VSS.n1130 VSS.n1129 585
R451 VSS.n4713 VSS.n1130 585
R452 VSS.n4715 VSS.n4714 585
R453 VSS.n4714 VSS.n4713 585
R454 VSS.n4709 VSS.n1198 585
R455 VSS.n4713 VSS.n1198 585
R456 VSS.n4712 VSS.n4711 585
R457 VSS.n4713 VSS.n4712 585
R458 VSS.n2681 VSS.n1131 585
R459 VSS.n1201 VSS.n1131 585
R460 VSS.n2844 VSS.n1131 585
R461 VSS.n1197 VSS.n1131 585
R462 VSS.n4766 VSS.n1131 585
R463 VSS.n4734 VSS.n1131 585
R464 VSS.n3267 VSS.n1131 585
R465 VSS.n3970 VSS.n1131 585
R466 VSS.n1836 VSS.n1131 585
R467 VSS.n4214 VSS.n1131 585
R468 VSS.n4709 VSS.n1208 585
R469 VSS.n4709 VSS.n4708 585
R470 VSS.n4716 VSS.n4715 585
R471 VSS.n4716 VSS.n1129 585
R472 VSS.n4718 VSS.n4715 585
R473 VSS.n4718 VSS.n1129 585
R474 VSS.n4719 VSS.n4718 585
R475 VSS.n4730 VSS.n1163 585
R476 VSS.n4730 VSS.n4729 585
R477 VSS.n4073 VSS.n3999 585
R478 VSS.n4073 VSS.n4072 585
R479 VSS.n5253 VSS.n298 585
R480 VSS.n302 VSS.n298 585
R481 VSS.n1227 VSS.n298 585
R482 VSS.n5046 VSS.n726 585
R483 VSS.n1306 VSS.n726 585
R484 VSS.n5013 VSS.n726 585
R485 VSS.n5009 VSS.n739 585
R486 VSS.n3870 VSS.n739 585
R487 VSS.n742 VSS.n739 585
R488 VSS.n4420 VSS.n1562 585
R489 VSS.n1566 VSS.n1562 585
R490 VSS.n4047 VSS.n1562 585
R491 VSS.n1566 VSS.n733 585
R492 VSS.n5011 VSS.n733 585
R493 VSS.n4420 VSS.n734 585
R494 VSS.n5011 VSS.n734 585
R495 VSS.n742 VSS.n732 585
R496 VSS.n5011 VSS.n732 585
R497 VSS.n5010 VSS.n5009 585
R498 VSS.n5011 VSS.n5010 585
R499 VSS.n5013 VSS.n5012 585
R500 VSS.n5012 VSS.n5011 585
R501 VSS.n5046 VSS.n724 585
R502 VSS.n5011 VSS.n724 585
R503 VSS.n698 VSS.n302 585
R504 VSS.n5011 VSS.n698 585
R505 VSS.n5253 VSS.n296 585
R506 VSS.n5011 VSS.n296 585
R507 VSS.n5287 VSS.n269 585
R508 VSS.n5255 VSS.n269 585
R509 VSS.n5080 VSS.n269 585
R510 VSS.n5048 VSS.n269 585
R511 VSS.n731 VSS.n269 585
R512 VSS.n735 VSS.n269 585
R513 VSS.n4454 VSS.n269 585
R514 VSS.n4422 VSS.n269 585
R515 VSS.n4319 VSS.n269 585
R516 VSS.n2514 VSS.n269 585
R517 VSS.n5253 VSS.n297 585
R518 VSS.n302 VSS.n297 585
R519 VSS.n5253 VSS.n5252 585
R520 VSS.n5252 VSS.n302 585
R521 VSS.n5252 VSS.n5251 585
R522 VSS.n5046 VSS.n725 585
R523 VSS.n5013 VSS.n725 585
R524 VSS.n5046 VSS.n5045 585
R525 VSS.n5045 VSS.n5013 585
R526 VSS.n5045 VSS.n5044 585
R527 VSS.n5009 VSS.n738 585
R528 VSS.n742 VSS.n738 585
R529 VSS.n5009 VSS.n5008 585
R530 VSS.n5008 VSS.n742 585
R531 VSS.n5008 VSS.n5007 585
R532 VSS.n4420 VSS.n1561 585
R533 VSS.n1566 VSS.n1561 585
R534 VSS.n4420 VSS.n4419 585
R535 VSS.n4419 VSS.n1566 585
R536 VSS.n4419 VSS.n4418 585
R537 VSS.n1389 VSS.n1387 585
R538 VSS.n1389 VSS.n209 585
R539 VSS.n4585 VSS.n1389 585
R540 VSS.n5535 VSS.n24 585
R541 VSS.n5535 VSS.n23 585
R542 VSS.n5536 VSS.n5535 585
R543 VSS.n5427 VSS.n5426 585
R544 VSS.n5428 VSS.n5427 585
R545 VSS.n5214 VSS.n5213 585
R546 VSS.n5215 VSS.n5214 585
R547 VSS.n4961 VSS.n4960 585
R548 VSS.n4962 VSS.n4961 585
R549 VSS.n5463 VSS.n57 585
R550 VSS.n5463 VSS.n13 585
R551 VSS.n5439 VSS.n13 585
R552 VSS.n5473 VSS.n57 585
R553 VSS.n5474 VSS.n5473 585
R554 VSS.n5473 VSS.n5472 585
R555 VSS.n4960 VSS.n4959 585
R556 VSS.n4959 VSS.n811 585
R557 VSS.n4959 VSS.n4958 585
R558 VSS.n5213 VSS.n5212 585
R559 VSS.n5212 VSS.n396 585
R560 VSS.n5212 VSS.n5211 585
R561 VSS.n5426 VSS.n5425 585
R562 VSS.n5425 VSS.n97 585
R563 VSS.n5425 VSS.n5424 585
R564 VSS.n5370 VSS.n5369 585
R565 VSS.n5373 VSS.n5372 585
R566 VSS.n5372 VSS.n5371 585
R567 VSS.n125 VSS.n123 585
R568 VSS.n127 VSS.n125 585
R569 VSS.n5411 VSS.n5410 585
R570 VSS.n5410 VSS.n5409 585
R571 VSS.n130 VSS.n126 585
R572 VSS.n5408 VSS.n126 585
R573 VSS.n5406 VSS.n5405 585
R574 VSS.n5407 VSS.n5406 585
R575 VSS.n133 VSS.n129 585
R576 VSS.n129 VSS.n128 585
R577 VSS.n5400 VSS.n5399 585
R578 VSS.n5399 VSS.n5398 585
R579 VSS.n5388 VSS.n134 585
R580 VSS.n5397 VSS.n134 585
R581 VSS.n5395 VSS.n5394 585
R582 VSS.n5396 VSS.n5395 585
R583 VSS.n5387 VSS.n102 585
R584 VSS.n5387 VSS.n5386 585
R585 VSS.n5418 VSS.n100 585
R586 VSS.n100 VSS.n99 585
R587 VSS.n5422 VSS.n5421 585
R588 VSS.n5423 VSS.n5422 585
R589 VSS.n5163 VSS.n96 585
R590 VSS.n5164 VSS.n5163 585
R591 VSS.n5161 VSS.n5159 585
R592 VSS.n5165 VSS.n5161 585
R593 VSS.n5198 VSS.n5197 585
R594 VSS.n5197 VSS.n5196 585
R595 VSS.n5168 VSS.n5162 585
R596 VSS.n5195 VSS.n5162 585
R597 VSS.n5193 VSS.n5192 585
R598 VSS.n5194 VSS.n5193 585
R599 VSS.n5171 VSS.n5167 585
R600 VSS.n5167 VSS.n5166 585
R601 VSS.n5187 VSS.n5186 585
R602 VSS.n5186 VSS.n5185 585
R603 VSS.n5175 VSS.n5172 585
R604 VSS.n5184 VSS.n5172 585
R605 VSS.n5182 VSS.n5181 585
R606 VSS.n5183 VSS.n5182 585
R607 VSS.n5174 VSS.n401 585
R608 VSS.n5174 VSS.n5173 585
R609 VSS.n5205 VSS.n399 585
R610 VSS.n399 VSS.n398 585
R611 VSS.n5209 VSS.n5208 585
R612 VSS.n5210 VSS.n5209 585
R613 VSS.n4910 VSS.n395 585
R614 VSS.n4911 VSS.n4910 585
R615 VSS.n4908 VSS.n4906 585
R616 VSS.n4912 VSS.n4908 585
R617 VSS.n4945 VSS.n4944 585
R618 VSS.n4944 VSS.n4943 585
R619 VSS.n4915 VSS.n4909 585
R620 VSS.n4942 VSS.n4909 585
R621 VSS.n4940 VSS.n4939 585
R622 VSS.n4941 VSS.n4940 585
R623 VSS.n4918 VSS.n4914 585
R624 VSS.n4914 VSS.n4913 585
R625 VSS.n4934 VSS.n4933 585
R626 VSS.n4933 VSS.n4932 585
R627 VSS.n4922 VSS.n4919 585
R628 VSS.n4931 VSS.n4919 585
R629 VSS.n4929 VSS.n4928 585
R630 VSS.n4930 VSS.n4929 585
R631 VSS.n4921 VSS.n816 585
R632 VSS.n4921 VSS.n4920 585
R633 VSS.n4952 VSS.n814 585
R634 VSS.n814 VSS.n813 585
R635 VSS.n4956 VSS.n4955 585
R636 VSS.n4957 VSS.n4956 585
R637 VSS.n3627 VSS.n810 585
R638 VSS.n3628 VSS.n3627 585
R639 VSS.n3625 VSS.n3623 585
R640 VSS.n3629 VSS.n3625 585
R641 VSS.n3667 VSS.n3666 585
R642 VSS.n3666 VSS.n3665 585
R643 VSS.n3632 VSS.n3626 585
R644 VSS.n3664 VSS.n3626 585
R645 VSS.n3662 VSS.n3661 585
R646 VSS.n3663 VSS.n3662 585
R647 VSS.n3635 VSS.n3631 585
R648 VSS.n3631 VSS.n3630 585
R649 VSS.n3656 VSS.n3655 585
R650 VSS.n3655 VSS.n3654 585
R651 VSS.n3639 VSS.n3636 585
R652 VSS.n3653 VSS.n3636 585
R653 VSS.n3651 VSS.n3650 585
R654 VSS.n3652 VSS.n3651 585
R655 VSS.n3644 VSS.n3638 585
R656 VSS.n3638 VSS.n3637 585
R657 VSS.n3645 VSS.n61 585
R658 VSS.n61 VSS.n60 585
R659 VSS.n5470 VSS.n5469 585
R660 VSS.n5471 VSS.n5470 585
R661 VSS.n5477 VSS.n5476 585
R662 VSS.n5476 VSS.n5475 585
R663 VSS.n5478 VSS.n52 585
R664 VSS.n52 VSS.n51 585
R665 VSS.n5490 VSS.n5489 585
R666 VSS.n5491 VSS.n5490 585
R667 VSS.n54 VSS.n48 585
R668 VSS.n5492 VSS.n48 585
R669 VSS.n5494 VSS.n50 585
R670 VSS.n5494 VSS.n5493 585
R671 VSS.n5495 VSS.n47 585
R672 VSS.n5495 VSS.n14 585
R673 VSS.n5497 VSS.n5496 585
R674 VSS.n5496 VSS.n15 585
R675 VSS.n44 VSS.n39 585
R676 VSS.n39 VSS.n38 585
R677 VSS.n5507 VSS.n5506 585
R678 VSS.n5508 VSS.n5507 585
R679 VSS.n41 VSS.n37 585
R680 VSS.n5509 VSS.n37 585
R681 VSS.n5512 VSS.n5511 585
R682 VSS.n5511 VSS.n5510 585
R683 VSS.n5513 VSS.n5 585
R684 VSS.n5 VSS.n3 585
R685 VSS.n2590 VSS.n2589 585
R686 VSS.n2620 VSS.n2619 585
R687 VSS.n2592 VSS.n2591 585
R688 VSS.n2618 VSS.n2592 585
R689 VSS.n2616 VSS.n2615 585
R690 VSS.n2617 VSS.n2616 585
R691 VSS.n2614 VSS.n2594 585
R692 VSS.n2594 VSS.n2593 585
R693 VSS.n2613 VSS.n2612 585
R694 VSS.n2612 VSS.n2611 585
R695 VSS.n2610 VSS.n2595 585
R696 VSS.n2610 VSS.n2609 585
R697 VSS.n2603 VSS.n2596 585
R698 VSS.n2608 VSS.n2596 585
R699 VSS.n2606 VSS.n2605 585
R700 VSS.n2607 VSS.n2606 585
R701 VSS.n2604 VSS.n2602 585
R702 VSS.n2602 VSS.n2597 585
R703 VSS.n2601 VSS.n2581 585
R704 VSS.n2601 VSS.n2600 585
R705 VSS.n2599 VSS.n2598 585
R706 VSS.n2677 VSS.n1858 585
R707 VSS.n2676 VSS.n1857 585
R708 VSS.n2580 VSS.n2579 585
R709 VSS.n2686 VSS.n2685 585
R710 VSS.n2687 VSS.n2686 585
R711 VSS.n2578 VSS.n2577 585
R712 VSS.n2688 VSS.n2578 585
R713 VSS.n2691 VSS.n2690 585
R714 VSS.n2690 VSS.n2689 585
R715 VSS.n2692 VSS.n2576 585
R716 VSS.n2576 VSS.n1181 585
R717 VSS.n2694 VSS.n2693 585
R718 VSS.n2694 VSS.n1180 585
R719 VSS.n2695 VSS.n2575 585
R720 VSS.n2696 VSS.n2695 585
R721 VSS.n2699 VSS.n2698 585
R722 VSS.n2698 VSS.n2697 585
R723 VSS.n2700 VSS.n2574 585
R724 VSS.n2574 VSS.n2573 585
R725 VSS.n2703 VSS.n2702 585
R726 VSS.n2704 VSS.n2703 585
R727 VSS.n2701 VSS.n2571 585
R728 VSS.n2705 VSS.n2571 585
R729 VSS.n2707 VSS.n2572 585
R730 VSS.n2707 VSS.n2706 585
R731 VSS.n2570 VSS.n2240 585
R732 VSS.n2570 VSS.n2569 585
R733 VSS.n2244 VSS.n2241 585
R734 VSS.n2568 VSS.n2241 585
R735 VSS.n2566 VSS.n2565 585
R736 VSS.n2567 VSS.n2566 585
R737 VSS.n2564 VSS.n2243 585
R738 VSS.n2243 VSS.n2242 585
R739 VSS.n2563 VSS.n2562 585
R740 VSS.n2562 VSS.n2561 585
R741 VSS.n2559 VSS.n2245 585
R742 VSS.n2560 VSS.n2559 585
R743 VSS.n2558 VSS.n2247 585
R744 VSS.n2558 VSS.n2557 585
R745 VSS.n2250 VSS.n2246 585
R746 VSS.n2556 VSS.n2246 585
R747 VSS.n2554 VSS.n2553 585
R748 VSS.n2555 VSS.n2554 585
R749 VSS.n2552 VSS.n2249 585
R750 VSS.n2249 VSS.n2248 585
R751 VSS.n2551 VSS.n2550 585
R752 VSS.n2550 VSS.n2549 585
R753 VSS.n2548 VSS.n2253 585
R754 VSS.n2547 VSS.n268 585
R755 VSS.n2389 VSS.n2388 585
R756 VSS.n2386 VSS.n2254 585
R757 VSS.n2385 VSS.n2256 585
R758 VSS.n2385 VSS.n2384 585
R759 VSS.n2259 VSS.n2255 585
R760 VSS.n2383 VSS.n2255 585
R761 VSS.n2381 VSS.n2380 585
R762 VSS.n2382 VSS.n2381 585
R763 VSS.n2379 VSS.n2258 585
R764 VSS.n2258 VSS.n2257 585
R765 VSS.n2378 VSS.n2377 585
R766 VSS.n2377 VSS.n2376 585
R767 VSS.n2261 VSS.n2260 585
R768 VSS.n2375 VSS.n2261 585
R769 VSS.n2373 VSS.n2372 585
R770 VSS.n2374 VSS.n2373 585
R771 VSS.n2371 VSS.n2263 585
R772 VSS.n2263 VSS.n2262 585
R773 VSS.n2370 VSS.n2369 585
R774 VSS.n2369 VSS.n2368 585
R775 VSS.n2367 VSS.n2366 585
R776 VSS.n2364 VSS.n1391 585
R777 VSS.n2265 VSS.n1390 585
R778 VSS.n2270 VSS.n2268 585
R779 VSS.n2322 VSS.n2321 585
R780 VSS.n2321 VSS.n2320 585
R781 VSS.n2269 VSS.n2266 585
R782 VSS.n2319 VSS.n2269 585
R783 VSS.n2317 VSS.n2316 585
R784 VSS.n2318 VSS.n2317 585
R785 VSS.n2315 VSS.n2272 585
R786 VSS.n2272 VSS.n2271 585
R787 VSS.n2314 VSS.n2313 585
R788 VSS.n2313 VSS.n2312 585
R789 VSS.n2274 VSS.n2273 585
R790 VSS.n2311 VSS.n2274 585
R791 VSS.n2309 VSS.n2308 585
R792 VSS.n2310 VSS.n2309 585
R793 VSS.n2307 VSS.n2276 585
R794 VSS.n2276 VSS.n2275 585
R795 VSS.n2306 VSS.n2305 585
R796 VSS.n2305 VSS.n2304 585
R797 VSS.n2303 VSS.n2278 585
R798 VSS.n2302 VSS.n2301 585
R799 VSS.n2286 VSS.n2279 585
R800 VSS.n2296 VSS.n2295 585
R801 VSS.n2289 VSS.n2285 585
R802 VSS.n2294 VSS.n2285 585
R803 VSS.n2292 VSS.n2291 585
R804 VSS.n2293 VSS.n2292 585
R805 VSS.n2290 VSS.n2288 585
R806 VSS.n2288 VSS.n2287 585
R807 VSS.n162 VSS.n160 585
R808 VSS.n160 VSS.n158 585
R809 VSS.n5384 VSS.n5383 585
R810 VSS.n5385 VSS.n5384 585
R811 VSS.n5382 VSS.n161 585
R812 VSS.n161 VSS.n159 585
R813 VSS.n5381 VSS.n5380 585
R814 VSS.n5380 VSS.n5379 585
R815 VSS.n164 VSS.n163 585
R816 VSS.n5378 VSS.n164 585
R817 VSS.n5376 VSS.n5375 585
R818 VSS.n5377 VSS.n5376 585
R819 VSS.n166 VSS.n165 585
R820 VSS.n4151 VSS.n1868 585
R821 VSS.n4152 VSS.n4151 585
R822 VSS.n4150 VSS.n4149 585
R823 VSS.n4150 VSS.n1900 585
R824 VSS.n4128 VSS.n1901 585
R825 VSS.n4122 VSS.n1901 585
R826 VSS.n4125 VSS.n4124 585
R827 VSS.n4124 VSS.n4123 585
R828 VSS.n4114 VSS.n1903 585
R829 VSS.n4121 VSS.n1903 585
R830 VSS.n4119 VSS.n4118 585
R831 VSS.n4120 VSS.n4119 585
R832 VSS.n1905 VSS.n1904 585
R833 VSS.n4106 VSS.n1904 585
R834 VSS.n4109 VSS.n4108 585
R835 VSS.n4108 VSS.n4107 585
R836 VSS.n4098 VSS.n1907 585
R837 VSS.n4105 VSS.n1907 585
R838 VSS.n4103 VSS.n4102 585
R839 VSS.n4104 VSS.n4103 585
R840 VSS.n1910 VSS.n1909 585
R841 VSS.n1909 VSS.n1908 585
R842 VSS.n4080 VSS.n4079 585
R843 VSS.n4079 VSS.n4078 585
R844 VSS.n3220 VSS.n1912 585
R845 VSS.n3222 VSS.n1912 585
R846 VSS.n3225 VSS.n3224 585
R847 VSS.n3224 VSS.n3223 585
R848 VSS.n3227 VSS.n3198 585
R849 VSS.n3198 VSS.n3197 585
R850 VSS.n3231 VSS.n3230 585
R851 VSS.n3232 VSS.n3231 585
R852 VSS.n3199 VSS.n3196 585
R853 VSS.n3233 VSS.n3196 585
R854 VSS.n3236 VSS.n3235 585
R855 VSS.n3235 VSS.n3234 585
R856 VSS.n3194 VSS.n3189 585
R857 VSS.n3189 VSS.n3188 585
R858 VSS.n3242 VSS.n3241 585
R859 VSS.n3243 VSS.n3242 585
R860 VSS.n3190 VSS.n1957 585
R861 VSS.n3244 VSS.n1957 585
R862 VSS.n3247 VSS.n3246 585
R863 VSS.n3246 VSS.n3245 585
R864 VSS.n1956 VSS.n1954 585
R865 VSS.n3187 VSS.n1956 585
R866 VSS.n3185 VSS.n3184 585
R867 VSS.n3186 VSS.n3185 585
R868 VSS.n3150 VSS.n3149 585
R869 VSS.n3149 VSS.n3148 585
R870 VSS.n3142 VSS.n1980 585
R871 VSS.n3147 VSS.n1980 585
R872 VSS.n3145 VSS.n3144 585
R873 VSS.n3146 VSS.n3145 585
R874 VSS.n3139 VSS.n1982 585
R875 VSS.n1982 VSS.n1981 585
R876 VSS.n1986 VSS.n1983 585
R877 VSS.n3131 VSS.n1986 585
R878 VSS.n3134 VSS.n3133 585
R879 VSS.n3133 VSS.n3132 585
R880 VSS.n3123 VSS.n1985 585
R881 VSS.n3130 VSS.n1985 585
R882 VSS.n3128 VSS.n3127 585
R883 VSS.n3129 VSS.n3128 585
R884 VSS.n1989 VSS.n1988 585
R885 VSS.n1988 VSS.n1987 585
R886 VSS.n3118 VSS.n3117 585
R887 VSS.n3117 VSS.n3116 585
R888 VSS.n3110 VSS.n1991 585
R889 VSS.n3115 VSS.n1991 585
R890 VSS.n3113 VSS.n3112 585
R891 VSS.n3114 VSS.n3113 585
R892 VSS.n3064 VSS.n3063 585
R893 VSS.n3063 VSS.n3062 585
R894 VSS.n2000 VSS.n1996 585
R895 VSS.n3061 VSS.n1996 585
R896 VSS.n3059 VSS.n3058 585
R897 VSS.n3060 VSS.n3059 585
R898 VSS.n2804 VSS.n1998 585
R899 VSS.n1998 VSS.n1997 585
R900 VSS.n2809 VSS.n2808 585
R901 VSS.n2810 VSS.n2809 585
R902 VSS.n2813 VSS.n2812 585
R903 VSS.n2812 VSS.n2811 585
R904 VSS.n2802 VSS.n2797 585
R905 VSS.n2797 VSS.n2796 585
R906 VSS.n2819 VSS.n2818 585
R907 VSS.n2820 VSS.n2819 585
R908 VSS.n2798 VSS.n2033 585
R909 VSS.n2821 VSS.n2033 585
R910 VSS.n2824 VSS.n2823 585
R911 VSS.n2823 VSS.n2822 585
R912 VSS.n2032 VSS.n2030 585
R913 VSS.n2795 VSS.n2032 585
R914 VSS.n2793 VSS.n2792 585
R915 VSS.n2794 VSS.n2793 585
R916 VSS.n2758 VSS.n2757 585
R917 VSS.n2757 VSS.n2756 585
R918 VSS.n2043 VSS.n2039 585
R919 VSS.n2755 VSS.n2039 585
R920 VSS.n2753 VSS.n2752 585
R921 VSS.n2754 VSS.n2753 585
R922 VSS.n2635 VSS.n2041 585
R923 VSS.n2041 VSS.n2040 585
R924 VSS.n2640 VSS.n2639 585
R925 VSS.n2641 VSS.n2640 585
R926 VSS.n2644 VSS.n2643 585
R927 VSS.n2643 VSS.n2642 585
R928 VSS.n2633 VSS.n2628 585
R929 VSS.n2628 VSS.n2627 585
R930 VSS.n2650 VSS.n2649 585
R931 VSS.n2651 VSS.n2650 585
R932 VSS.n2629 VSS.n2588 585
R933 VSS.n2652 VSS.n2588 585
R934 VSS.n2655 VSS.n2654 585
R935 VSS.n2654 VSS.n2653 585
R936 VSS.n2587 VSS.n2585 585
R937 VSS.n2626 VSS.n2587 585
R938 VSS.n2624 VSS.n2623 585
R939 VSS.n2625 VSS.n2624 585
R940 VSS.n4157 VSS.n4156 585
R941 VSS.n4154 VSS.n1869 585
R942 VSS.n4178 VSS.n4177 585
R943 VSS.n4176 VSS.n1853 585
R944 VSS.n4176 VSS.n1859 585
R945 VSS.n4175 VSS.n1861 585
R946 VSS.n4175 VSS.n4174 585
R947 VSS.n4169 VSS.n1860 585
R948 VSS.n4173 VSS.n1860 585
R949 VSS.n4171 VSS.n4170 585
R950 VSS.n4172 VSS.n4171 585
R951 VSS.n4168 VSS.n1863 585
R952 VSS.n1863 VSS.n1862 585
R953 VSS.n4167 VSS.n4166 585
R954 VSS.n4166 VSS.n4165 585
R955 VSS.n1865 VSS.n1864 585
R956 VSS.n4164 VSS.n1865 585
R957 VSS.n4162 VSS.n4161 585
R958 VSS.n4163 VSS.n4162 585
R959 VSS.n4160 VSS.n1867 585
R960 VSS.n1867 VSS.n1866 585
R961 VSS.n4179 VSS.n1850 585
R962 VSS.n4193 VSS.n4192 585
R963 VSS.n4192 VSS.n4191 585
R964 VSS.n4194 VSS.n4188 585
R965 VSS.n4188 VSS.n4187 585
R966 VSS.n4196 VSS.n4195 585
R967 VSS.n4197 VSS.n4196 585
R968 VSS.n4189 VSS.n4186 585
R969 VSS.n4198 VSS.n4186 585
R970 VSS.n4200 VSS.n4185 585
R971 VSS.n4200 VSS.n4199 585
R972 VSS.n4202 VSS.n4201 585
R973 VSS.n4201 VSS.n1184 585
R974 VSS.n4203 VSS.n4184 585
R975 VSS.n4184 VSS.n1183 585
R976 VSS.n4205 VSS.n4204 585
R977 VSS.n4206 VSS.n4205 585
R978 VSS.n1856 VSS.n1854 585
R979 VSS.n4207 VSS.n1856 585
R980 VSS.n4210 VSS.n4209 585
R981 VSS.n4209 VSS.n4208 585
R982 VSS.n4183 VSS.n1855 585
R983 VSS.n4182 VSS.n4181 585
R984 VSS.n4190 VSS.n1359 585
R985 VSS.n1359 VSS.n1358 585
R986 VSS.n2527 VSS.n2521 585
R987 VSS.n2530 VSS.n2529 585
R988 VSS.n2529 VSS.n2528 585
R989 VSS.n2519 VSS.n2518 585
R990 VSS.n2526 VSS.n2519 585
R991 VSS.n2524 VSS.n2523 585
R992 VSS.n2525 VSS.n2524 585
R993 VSS.n2522 VSS.n1366 585
R994 VSS.n1368 VSS.n1366 585
R995 VSS.n4666 VSS.n1367 585
R996 VSS.n4666 VSS.n4665 585
R997 VSS.n4667 VSS.n1365 585
R998 VSS.n4668 VSS.n4667 585
R999 VSS.n4671 VSS.n4670 585
R1000 VSS.n4670 VSS.n4669 585
R1001 VSS.n4672 VSS.n1364 585
R1002 VSS.n1364 VSS.n1363 585
R1003 VSS.n4674 VSS.n4673 585
R1004 VSS.n4675 VSS.n4674 585
R1005 VSS.n1362 VSS.n1361 585
R1006 VSS.n4676 VSS.n1362 585
R1007 VSS.n4679 VSS.n4678 585
R1008 VSS.n4678 VSS.n4677 585
R1009 VSS.n2392 VSS.n2390 585
R1010 VSS.n4645 VSS.n1386 585
R1011 VSS.n1386 VSS.n1385 585
R1012 VSS.n4647 VSS.n4646 585
R1013 VSS.n4648 VSS.n4647 585
R1014 VSS.n1384 VSS.n1383 585
R1015 VSS.n4649 VSS.n1384 585
R1016 VSS.n4652 VSS.n4651 585
R1017 VSS.n4651 VSS.n4650 585
R1018 VSS.n4653 VSS.n1381 585
R1019 VSS.n1381 VSS.n1379 585
R1020 VSS.n4655 VSS.n4654 585
R1021 VSS.n4656 VSS.n4655 585
R1022 VSS.n1382 VSS.n1380 585
R1023 VSS.n2533 VSS.n1380 585
R1024 VSS.n2536 VSS.n2535 585
R1025 VSS.n2537 VSS.n2536 585
R1026 VSS.n2534 VSS.n2517 585
R1027 VSS.n2538 VSS.n2517 585
R1028 VSS.n2540 VSS.n2532 585
R1029 VSS.n2540 VSS.n2539 585
R1030 VSS.n2541 VSS.n2391 585
R1031 VSS.n2544 VSS.n2543 585
R1032 VSS.n4644 VSS.n4643 585
R1033 VSS.n4643 VSS.n4642 585
R1034 VSS.n4597 VSS.n4596 585
R1035 VSS.n4599 VSS.n4597 585
R1036 VSS.n4602 VSS.n4601 585
R1037 VSS.n4601 VSS.n4600 585
R1038 VSS.n4603 VSS.n4593 585
R1039 VSS.n4593 VSS.n4592 585
R1040 VSS.n4605 VSS.n4604 585
R1041 VSS.n4606 VSS.n4605 585
R1042 VSS.n4594 VSS.n4591 585
R1043 VSS.n4607 VSS.n4591 585
R1044 VSS.n4609 VSS.n4590 585
R1045 VSS.n4609 VSS.n4608 585
R1046 VSS.n4612 VSS.n4611 585
R1047 VSS.n4611 VSS.n4610 585
R1048 VSS.n4613 VSS.n1406 585
R1049 VSS.n1406 VSS.n1404 585
R1050 VSS.n4615 VSS.n4614 585
R1051 VSS.n4616 VSS.n4615 585
R1052 VSS.n4589 VSS.n1405 585
R1053 VSS.n1405 VSS.n1403 585
R1054 VSS.n4588 VSS.n4587 585
R1055 VSS.n4587 VSS.n1392 585
R1056 VSS.n4586 VSS.n1388 585
R1057 VSS.n4640 VSS.n1388 585
R1058 VSS.n4595 VSS.n21 585
R1059 VSS.n4598 VSS.n21 585
R1060 VSS.n5560 VSS.n4 585
R1061 VSS.n5559 VSS.n8 585
R1062 VSS.n5559 VSS.n5558 585
R1063 VSS.n5553 VSS.n7 585
R1064 VSS.n5557 VSS.n7 585
R1065 VSS.n5555 VSS.n5554 585
R1066 VSS.n5556 VSS.n5555 585
R1067 VSS.n5552 VSS.n10 585
R1068 VSS.n10 VSS.n9 585
R1069 VSS.n5551 VSS.n5550 585
R1070 VSS.n5550 VSS.n5549 585
R1071 VSS.n12 VSS.n11 585
R1072 VSS.n5548 VSS.n12 585
R1073 VSS.n5546 VSS.n5545 585
R1074 VSS.n5547 VSS.n5546 585
R1075 VSS.n5544 VSS.n17 585
R1076 VSS.n17 VSS.n16 585
R1077 VSS.n5543 VSS.n5542 585
R1078 VSS.n5542 VSS.n5541 585
R1079 VSS.n19 VSS.n18 585
R1080 VSS.n5540 VSS.n19 585
R1081 VSS.n5538 VSS.n5537 585
R1082 VSS.n5539 VSS.n5538 585
R1083 VSS.n5563 VSS.n5562 585
R1084 VSS.n2619 VSS.n2589 578.947
R1085 VSS.n2619 VSS.n2618 578.947
R1086 VSS.n2618 VSS.n2617 578.947
R1087 VSS.n2617 VSS.n2593 578.947
R1088 VSS.n2611 VSS.n2593 578.947
R1089 VSS.n2609 VSS.n2608 578.947
R1090 VSS.n2608 VSS.n2607 578.947
R1091 VSS.n2607 VSS.n2597 578.947
R1092 VSS.n2600 VSS.n2597 578.947
R1093 VSS.n2600 VSS.n2599 578.947
R1094 VSS.n2599 VSS.n1858 578.947
R1095 VSS.n2579 VSS.n1857 578.947
R1096 VSS.n2687 VSS.n2579 578.947
R1097 VSS.n2688 VSS.n2687 578.947
R1098 VSS.n2689 VSS.n2688 578.947
R1099 VSS.n2689 VSS.n1181 578.947
R1100 VSS.n2696 VSS.n1180 578.947
R1101 VSS.n2697 VSS.n2696 578.947
R1102 VSS.n2697 VSS.n2573 578.947
R1103 VSS.n2704 VSS.n2573 578.947
R1104 VSS.n2705 VSS.n2704 578.947
R1105 VSS.n2706 VSS.n2705 578.947
R1106 VSS.n2569 VSS.n2568 578.947
R1107 VSS.n2568 VSS.n2567 578.947
R1108 VSS.n2567 VSS.n2242 578.947
R1109 VSS.n2561 VSS.n2242 578.947
R1110 VSS.n2561 VSS.n2560 578.947
R1111 VSS.n2557 VSS.n2556 578.947
R1112 VSS.n2556 VSS.n2555 578.947
R1113 VSS.n2555 VSS.n2248 578.947
R1114 VSS.n2549 VSS.n2248 578.947
R1115 VSS.n2549 VSS.n2548 578.947
R1116 VSS.n2548 VSS.n2547 578.947
R1117 VSS.n2389 VSS.n2254 578.947
R1118 VSS.n2384 VSS.n2254 578.947
R1119 VSS.n2384 VSS.n2383 578.947
R1120 VSS.n2383 VSS.n2382 578.947
R1121 VSS.n2382 VSS.n2257 578.947
R1122 VSS.n2376 VSS.n2375 578.947
R1123 VSS.n2375 VSS.n2374 578.947
R1124 VSS.n2374 VSS.n2262 578.947
R1125 VSS.n2368 VSS.n2262 578.947
R1126 VSS.n2368 VSS.n2367 578.947
R1127 VSS.n2367 VSS.n1391 578.947
R1128 VSS.n2270 VSS.n1390 578.947
R1129 VSS.n2320 VSS.n2270 578.947
R1130 VSS.n2320 VSS.n2319 578.947
R1131 VSS.n2319 VSS.n2318 578.947
R1132 VSS.n2318 VSS.n2271 578.947
R1133 VSS.n2312 VSS.n2311 578.947
R1134 VSS.n2311 VSS.n2310 578.947
R1135 VSS.n2310 VSS.n2275 578.947
R1136 VSS.n2304 VSS.n2275 578.947
R1137 VSS.n2304 VSS.n2303 578.947
R1138 VSS.n2303 VSS.n2302 578.947
R1139 VSS.n2295 VSS.n2286 578.947
R1140 VSS.n2295 VSS.n2294 578.947
R1141 VSS.n2294 VSS.n2293 578.947
R1142 VSS.n2293 VSS.n2287 578.947
R1143 VSS.n2287 VSS.n158 578.947
R1144 VSS.n5385 VSS.n159 578.947
R1145 VSS.n5379 VSS.n159 578.947
R1146 VSS.n5379 VSS.n5378 578.947
R1147 VSS.n5378 VSS.n5377 578.947
R1148 VSS.n5377 VSS.n165 578.947
R1149 VSS.n1874 VSS.n1873 557.503
R1150 VSS.n4155 VSS.n1866 530.74
R1151 VSS.t83 VSS.n1890 517.26
R1152 VSS.n2777 VSS.t38 502.363
R1153 VSS.t33 VSS.n1173 502.363
R1154 VSS.t33 VSS.n1175 502.363
R1155 VSS.n1673 VSS.t44 502.363
R1156 VSS.n4975 VSS.t44 502.363
R1157 VSS.n664 VSS.t44 502.363
R1158 VSS.t33 VSS.n1178 502.363
R1159 VSS.n1862 VSS.t38 496.498
R1160 VSS.t33 VSS.n1184 496.498
R1161 VSS.n4180 VSS.n1858 482.457
R1162 VSS.n2706 VSS.n1265 482.457
R1163 VSS.n4641 VSS.n1391 482.457
R1164 VSS.n2302 VSS.n20 482.457
R1165 VSS.n5424 VSS.n5423 475.803
R1166 VSS.n5211 VSS.n5210 475.803
R1167 VSS.n4958 VSS.n4957 475.803
R1168 VSS.n5472 VSS.n5471 475.803
R1169 VSS.n4156 VSS.n4155 471.144
R1170 VSS.n4661 VSS.n4660 454.401
R1171 VSS.n4621 VSS.n1400 454.401
R1172 VSS.n5371 VSS.n5370 452.248
R1173 VSS.n5164 VSS.n97 452.248
R1174 VSS.n4911 VSS.n396 452.248
R1175 VSS.n3628 VSS.n811 452.248
R1176 VSS.n5475 VSS.n5474 452.248
R1177 VSS.t67 VSS.n1881 446.87
R1178 VSS.n5371 VSS.n127 423.983
R1179 VSS.n5409 VSS.n127 423.983
R1180 VSS.n5409 VSS.n5408 423.983
R1181 VSS.n5408 VSS.n5407 423.983
R1182 VSS.n5407 VSS.n128 423.983
R1183 VSS.n5398 VSS.n5397 423.983
R1184 VSS.n5397 VSS.n5396 423.983
R1185 VSS.n5396 VSS.n5386 423.983
R1186 VSS.n5386 VSS.n99 423.983
R1187 VSS.n5423 VSS.n99 423.983
R1188 VSS.n5165 VSS.n5164 423.983
R1189 VSS.n5196 VSS.n5165 423.983
R1190 VSS.n5196 VSS.n5195 423.983
R1191 VSS.n5195 VSS.n5194 423.983
R1192 VSS.n5194 VSS.n5166 423.983
R1193 VSS.n5185 VSS.n5184 423.983
R1194 VSS.n5184 VSS.n5183 423.983
R1195 VSS.n5183 VSS.n5173 423.983
R1196 VSS.n5173 VSS.n398 423.983
R1197 VSS.n5210 VSS.n398 423.983
R1198 VSS.n4912 VSS.n4911 423.983
R1199 VSS.n4943 VSS.n4912 423.983
R1200 VSS.n4943 VSS.n4942 423.983
R1201 VSS.n4942 VSS.n4941 423.983
R1202 VSS.n4941 VSS.n4913 423.983
R1203 VSS.n4932 VSS.n4931 423.983
R1204 VSS.n4931 VSS.n4930 423.983
R1205 VSS.n4930 VSS.n4920 423.983
R1206 VSS.n4920 VSS.n813 423.983
R1207 VSS.n4957 VSS.n813 423.983
R1208 VSS.n3629 VSS.n3628 423.983
R1209 VSS.n3665 VSS.n3629 423.983
R1210 VSS.n3665 VSS.n3664 423.983
R1211 VSS.n3664 VSS.n3663 423.983
R1212 VSS.n3663 VSS.n3630 423.983
R1213 VSS.n3654 VSS.n3653 423.983
R1214 VSS.n3653 VSS.n3652 423.983
R1215 VSS.n3652 VSS.n3637 423.983
R1216 VSS.n3637 VSS.n60 423.983
R1217 VSS.n5471 VSS.n60 423.983
R1218 VSS.n5475 VSS.n51 423.983
R1219 VSS.n5491 VSS.n51 423.983
R1220 VSS.n5492 VSS.n5491 423.983
R1221 VSS.n5493 VSS.n5492 423.983
R1222 VSS.n5493 VSS.n14 423.983
R1223 VSS.n38 VSS.n15 423.983
R1224 VSS.n5508 VSS.n38 423.983
R1225 VSS.n5509 VSS.n5508 423.983
R1226 VSS.n5510 VSS.n5509 423.983
R1227 VSS.n5510 VSS.n3 423.983
R1228 VSS.n1883 VSS.t82 414.101
R1229 VSS.n2626 VSS.n2625 396.795
R1230 VSS.n2653 VSS.n2626 396.795
R1231 VSS.n2653 VSS.n2652 396.795
R1232 VSS.n2652 VSS.n2651 396.795
R1233 VSS.n2651 VSS.n2627 396.795
R1234 VSS.n2642 VSS.n2641 396.795
R1235 VSS.n2641 VSS.n2040 396.795
R1236 VSS.n2754 VSS.n2040 396.795
R1237 VSS.n2755 VSS.n2754 396.795
R1238 VSS.n2756 VSS.n2755 396.795
R1239 VSS.n2795 VSS.n2794 396.795
R1240 VSS.n2822 VSS.n2795 396.795
R1241 VSS.n2822 VSS.n2821 396.795
R1242 VSS.n2821 VSS.n2820 396.795
R1243 VSS.n2820 VSS.n2796 396.795
R1244 VSS.n2811 VSS.n2810 396.795
R1245 VSS.n2810 VSS.n1997 396.795
R1246 VSS.n3060 VSS.n1997 396.795
R1247 VSS.n3061 VSS.n3060 396.795
R1248 VSS.n3062 VSS.n3061 396.795
R1249 VSS.n3115 VSS.n3114 396.795
R1250 VSS.n3116 VSS.n3115 396.795
R1251 VSS.n3116 VSS.n1987 396.795
R1252 VSS.n3129 VSS.n1987 396.795
R1253 VSS.n3130 VSS.n3129 396.795
R1254 VSS.n3132 VSS.n3131 396.795
R1255 VSS.n3131 VSS.n1981 396.795
R1256 VSS.n3146 VSS.n1981 396.795
R1257 VSS.n3147 VSS.n3146 396.795
R1258 VSS.n3148 VSS.n3147 396.795
R1259 VSS.n3187 VSS.n3186 396.795
R1260 VSS.n3245 VSS.n3187 396.795
R1261 VSS.n3245 VSS.n3244 396.795
R1262 VSS.n3244 VSS.n3243 396.795
R1263 VSS.n3243 VSS.n3188 396.795
R1264 VSS.n3234 VSS.n3233 396.795
R1265 VSS.n3233 VSS.n3232 396.795
R1266 VSS.n3232 VSS.n3197 396.795
R1267 VSS.n3223 VSS.n3197 396.795
R1268 VSS.n3223 VSS.n3222 396.795
R1269 VSS.n4078 VSS.n1908 396.795
R1270 VSS.n4104 VSS.n1908 396.795
R1271 VSS.n4105 VSS.n4104 396.795
R1272 VSS.n4107 VSS.n4105 396.795
R1273 VSS.n4107 VSS.n4106 396.795
R1274 VSS.n4121 VSS.n4120 396.795
R1275 VSS.n4123 VSS.n4121 396.795
R1276 VSS.n4123 VSS.n4122 396.795
R1277 VSS.n4122 VSS.n1900 396.795
R1278 VSS.n4152 VSS.n1900 396.795
R1279 VSS.n2611 VSS.t38 392.399
R1280 VSS.t33 VSS.n1181 392.399
R1281 VSS.n2560 VSS.t31 392.399
R1282 VSS.n2257 VSS.t40 392.399
R1283 VSS.n2271 VSS.t44 392.399
R1284 VSS.t42 VSS.n158 392.399
R1285 VSS.n1896 VSS.n1891 377.519
R1286 VSS.t42 VSS.n157 129
R1287 VSS.n803 VSS.t42 129
R1288 VSS.n388 VSS.t42 129
R1289 VSS.n5462 VSS.t42 129
R1290 VSS.n4659 VSS.n1377 326.163
R1291 VSS.n4662 VSS.n1371 325.788
R1292 VSS.n5428 VSS.t42 129.871
R1293 VSS.n4962 VSS.t42 129.871
R1294 VSS.n5215 VSS.t42 129.871
R1295 VSS.t42 VSS.n13 129.871
R1296 VSS.n4624 VSS.n4623 311.416
R1297 VSS.n5228 VSS.n334 292.5
R1298 VSS.n5221 VSS.n5220 292.5
R1299 VSS.n5223 VSS.n343 292.5
R1300 VSS.n354 VSS.n342 292.5
R1301 VSS.n356 VSS.n355 292.5
R1302 VSS.n353 VSS.n346 292.5
R1303 VSS.n352 VSS.n351 292.5
R1304 VSS.n350 VSS.n349 292.5
R1305 VSS.n348 VSS.n347 292.5
R1306 VSS.n337 VSS.n335 292.5
R1307 VSS.n5227 VSS.n5226 292.5
R1308 VSS.n5219 VSS.n5218 292.5
R1309 VSS.n393 VSS.n392 292.5
R1310 VSS.n391 VSS.n390 292.5
R1311 VSS.n370 VSS.n369 292.5
R1312 VSS.n386 VSS.n385 292.5
R1313 VSS.n384 VSS.n373 292.5
R1314 VSS.n383 VSS.n382 292.5
R1315 VSS.n381 VSS.n380 292.5
R1316 VSS.n379 VSS.n378 292.5
R1317 VSS.n377 VSS.n376 292.5
R1318 VSS.n375 VSS.n374 292.5
R1319 VSS.n5216 VSS.n361 292.5
R1320 VSS.n808 VSS.n807 292.5
R1321 VSS.n806 VSS.n805 292.5
R1322 VSS.n785 VSS.n784 292.5
R1323 VSS.n801 VSS.n800 292.5
R1324 VSS.n799 VSS.n788 292.5
R1325 VSS.n798 VSS.n797 292.5
R1326 VSS.n796 VSS.n795 292.5
R1327 VSS.n794 VSS.n793 292.5
R1328 VSS.n792 VSS.n791 292.5
R1329 VSS.n790 VSS.n789 292.5
R1330 VSS.n4963 VSS.n776 292.5
R1331 VSS.n4965 VSS.n774 292.5
R1332 VSS.n4966 VSS.n4965 292.5
R1333 VSS.n4969 VSS.n4968 292.5
R1334 VSS.n4968 VSS.n4967 292.5
R1335 VSS.n4970 VSS.n772 292.5
R1336 VSS.n772 VSS.n771 292.5
R1337 VSS.n4972 VSS.n4971 292.5
R1338 VSS.n4973 VSS.n4972 292.5
R1339 VSS.n773 VSS.n769 292.5
R1340 VSS.n4974 VSS.n769 292.5
R1341 VSS.n4976 VSS.n770 292.5
R1342 VSS.n4976 VSS.n4975 292.5
R1343 VSS.n4977 VSS.n768 292.5
R1344 VSS.n4978 VSS.n4977 292.5
R1345 VSS.n4981 VSS.n4980 292.5
R1346 VSS.n4980 VSS.n4979 292.5
R1347 VSS.n4982 VSS.n767 292.5
R1348 VSS.n767 VSS.n766 292.5
R1349 VSS.n4984 VSS.n4983 292.5
R1350 VSS.n4985 VSS.n4984 292.5
R1351 VSS.n765 VSS.n763 292.5
R1352 VSS.n4988 VSS.n4987 292.5
R1353 VSS.n2363 VSS.n2358 292.5
R1354 VSS.n1732 VSS.n1407 292.5
R1355 VSS.n1735 VSS.n1734 292.5
R1356 VSS.n1729 VSS.n1728 292.5
R1357 VSS.n1714 VSS.n1713 292.5
R1358 VSS.n1717 VSS.n1716 292.5
R1359 VSS.n4370 VSS.n4369 292.5
R1360 VSS.n4372 VSS.n1699 292.5
R1361 VSS.n4375 VSS.n4374 292.5
R1362 VSS.n1697 VSS.n1690 292.5
R1363 VSS.n4399 VSS.n4398 292.5
R1364 VSS.n1649 VSS.n1648 292.5
R1365 VSS.n1645 VSS.n1644 292.5
R1366 VSS.n1639 VSS.n1638 292.5
R1367 VSS.n1636 VSS.n1635 292.5
R1368 VSS.n1630 VSS.n1629 292.5
R1369 VSS.n1627 VSS.n1489 292.5
R1370 VSS.n4486 VSS.n4485 292.5
R1371 VSS.n4489 VSS.n4488 292.5
R1372 VSS.n1484 VSS.n1476 292.5
R1373 VSS.n1482 VSS.n1475 292.5
R1374 VSS.n3735 VSS.n3734 292.5
R1375 VSS.n3731 VSS.n3730 292.5
R1376 VSS.n3725 VSS.n3724 292.5
R1377 VSS.n3722 VSS.n3721 292.5
R1378 VSS.n3716 VSS.n3715 292.5
R1379 VSS.n3713 VSS.n1010 292.5
R1380 VSS.n4859 VSS.n4858 292.5
R1381 VSS.n4862 VSS.n4861 292.5
R1382 VSS.n1005 VSS.n997 292.5
R1383 VSS.n1003 VSS.n996 292.5
R1384 VSS.n940 VSS.n939 292.5
R1385 VSS.n936 VSS.n935 292.5
R1386 VSS.n930 VSS.n929 292.5
R1387 VSS.n927 VSS.n926 292.5
R1388 VSS.n921 VSS.n920 292.5
R1389 VSS.n918 VSS.n469 292.5
R1390 VSS.n5112 VSS.n5111 292.5
R1391 VSS.n5115 VSS.n5114 292.5
R1392 VSS.n639 VSS.n459 292.5
R1393 VSS.n641 VSS.n458 292.5
R1394 VSS.n637 VSS.n636 292.5
R1395 VSS.n633 VSS.n632 292.5
R1396 VSS.n622 VSS.n621 292.5
R1397 VSS.n619 VSS.n218 292.5
R1398 VSS.n617 VSS.n616 292.5
R1399 VSS.n5319 VSS.n5318 292.5
R1400 VSS.n5321 VSS.n210 292.5
R1401 VSS.n5324 VSS.n5323 292.5
R1402 VSS.n2359 VSS.n203 292.5
R1403 VSS.n2361 VSS.n202 292.5
R1404 VSS.n1663 VSS.n71 292.5
R1405 VSS.n1664 VSS.n71 292.5
R1406 VSS.n1667 VSS.n1666 292.5
R1407 VSS.n1666 VSS.n1665 292.5
R1408 VSS.n1668 VSS.n1661 292.5
R1409 VSS.n1661 VSS.n1660 292.5
R1410 VSS.n1670 VSS.n1669 292.5
R1411 VSS.n1671 VSS.n1670 292.5
R1412 VSS.n1662 VSS.n1658 292.5
R1413 VSS.n1672 VSS.n1658 292.5
R1414 VSS.n1674 VSS.n1659 292.5
R1415 VSS.n1674 VSS.n1673 292.5
R1416 VSS.n1675 VSS.n1657 292.5
R1417 VSS.n1676 VSS.n1675 292.5
R1418 VSS.n1679 VSS.n1678 292.5
R1419 VSS.n1678 VSS.n1677 292.5
R1420 VSS.n1680 VSS.n1656 292.5
R1421 VSS.n1656 VSS.n1655 292.5
R1422 VSS.n1682 VSS.n1681 292.5
R1423 VSS.n1683 VSS.n1682 292.5
R1424 VSS.n1654 VSS.n1652 292.5
R1425 VSS.n1686 VSS.n1685 292.5
R1426 VSS.n5533 VSS.n5532 292.5
R1427 VSS.n4548 VSS.n4547 292.5
R1428 VSS.n4545 VSS.n4543 292.5
R1429 VSS.n4558 VSS.n4557 292.5
R1430 VSS.n4560 VSS.n4533 292.5
R1431 VSS.n4563 VSS.n4562 292.5
R1432 VSS.n4531 VSS.n4529 292.5
R1433 VSS.n4573 VSS.n4572 292.5
R1434 VSS.n4576 VSS.n4575 292.5
R1435 VSS.n4505 VSS.n4504 292.5
R1436 VSS.n3542 VSS.n1453 292.5
R1437 VSS.n3545 VSS.n3544 292.5
R1438 VSS.n3550 VSS.n3549 292.5
R1439 VSS.n3552 VSS.n3517 292.5
R1440 VSS.n3555 VSS.n3554 292.5
R1441 VSS.n3533 VSS.n3532 292.5
R1442 VSS.n3527 VSS.n3526 292.5
R1443 VSS.n3524 VSS.n3523 292.5
R1444 VSS.n3675 VSS.n3674 292.5
R1445 VSS.n3677 VSS.n3479 292.5
R1446 VSS.n3684 VSS.n3683 292.5
R1447 VSS.n3474 VSS.n3473 292.5
R1448 VSS.n3468 VSS.n3467 292.5
R1449 VSS.n3465 VSS.n3464 292.5
R1450 VSS.n3459 VSS.n3458 292.5
R1451 VSS.n3456 VSS.n976 292.5
R1452 VSS.n4878 VSS.n4877 292.5
R1453 VSS.n4881 VSS.n4880 292.5
R1454 VSS.n971 VSS.n839 292.5
R1455 VSS.n969 VSS.n838 292.5
R1456 VSS.n963 VSS.n962 292.5
R1457 VSS.n872 VSS.n871 292.5
R1458 VSS.n869 VSS.n868 292.5
R1459 VSS.n854 VSS.n851 292.5
R1460 VSS.n857 VSS.n856 292.5
R1461 VSS.n852 VSS.n438 292.5
R1462 VSS.n5131 VSS.n5130 292.5
R1463 VSS.n5134 VSS.n5133 292.5
R1464 VSS.n433 VSS.n424 292.5
R1465 VSS.n431 VSS.n423 292.5
R1466 VSS.n594 VSS.n593 292.5
R1467 VSS.n590 VSS.n589 292.5
R1468 VSS.n584 VSS.n583 292.5
R1469 VSS.n581 VSS.n580 292.5
R1470 VSS.n575 VSS.n574 292.5
R1471 VSS.n5339 VSS.n5338 292.5
R1472 VSS.n5341 VSS.n178 292.5
R1473 VSS.n5344 VSS.n5343 292.5
R1474 VSS.n2280 VSS.n170 292.5
R1475 VSS.n2282 VSS.n169 292.5
R1476 VSS.n2298 VSS.n2284 292.5
R1477 VSS.n153 VSS.n152 292.5
R1478 VSS.n155 VSS.n154 292.5
R1479 VSS.n151 VSS.n138 292.5
R1480 VSS.n150 VSS.n149 292.5
R1481 VSS.n148 VSS.n147 292.5
R1482 VSS.n146 VSS.n145 292.5
R1483 VSS.n144 VSS.n143 292.5
R1484 VSS.n142 VSS.n141 292.5
R1485 VSS.n140 VSS.n139 292.5
R1486 VSS.n654 VSS.n82 292.5
R1487 VSS.n655 VSS.n654 292.5
R1488 VSS.n87 VSS.n85 292.5
R1489 VSS.n5430 VSS.n5429 292.5
R1490 VSS.n658 VSS.n657 292.5
R1491 VSS.n657 VSS.n656 292.5
R1492 VSS.n659 VSS.n652 292.5
R1493 VSS.n652 VSS.n651 292.5
R1494 VSS.n661 VSS.n660 292.5
R1495 VSS.n662 VSS.n661 292.5
R1496 VSS.n653 VSS.n649 292.5
R1497 VSS.n663 VSS.n649 292.5
R1498 VSS.n665 VSS.n650 292.5
R1499 VSS.n665 VSS.n664 292.5
R1500 VSS.n666 VSS.n648 292.5
R1501 VSS.n667 VSS.n666 292.5
R1502 VSS.n670 VSS.n669 292.5
R1503 VSS.n669 VSS.n668 292.5
R1504 VSS.n671 VSS.n647 292.5
R1505 VSS.n647 VSS.n646 292.5
R1506 VSS.n673 VSS.n672 292.5
R1507 VSS.n674 VSS.n673 292.5
R1508 VSS.n645 VSS.n644 292.5
R1509 VSS.n677 VSS.n676 292.5
R1510 VSS.n5237 VSS.n303 292.5
R1511 VSS.n5239 VSS.n5238 292.5
R1512 VSS.n319 VSS.n318 292.5
R1513 VSS.n317 VSS.n316 292.5
R1514 VSS.n315 VSS.n314 292.5
R1515 VSS.n313 VSS.n312 292.5
R1516 VSS.n5242 VSS.n309 292.5
R1517 VSS.n5245 VSS.n5244 292.5
R1518 VSS.n5247 VSS.n5246 292.5
R1519 VSS.n5249 VSS.n5248 292.5
R1520 VSS.n4993 VSS.n743 292.5
R1521 VSS.n4995 VSS.n4994 292.5
R1522 VSS.n759 VSS.n758 292.5
R1523 VSS.n757 VSS.n756 292.5
R1524 VSS.n755 VSS.n754 292.5
R1525 VSS.n753 VSS.n752 292.5
R1526 VSS.n4998 VSS.n749 292.5
R1527 VSS.n5001 VSS.n5000 292.5
R1528 VSS.n5003 VSS.n5002 292.5
R1529 VSS.n5005 VSS.n5004 292.5
R1530 VSS.n4404 VSS.n1567 292.5
R1531 VSS.n4406 VSS.n4405 292.5
R1532 VSS.n1583 VSS.n1582 292.5
R1533 VSS.n1581 VSS.n1580 292.5
R1534 VSS.n1579 VSS.n1578 292.5
R1535 VSS.n1577 VSS.n1576 292.5
R1536 VSS.n4409 VSS.n1573 292.5
R1537 VSS.n4412 VSS.n4411 292.5
R1538 VSS.n4414 VSS.n4413 292.5
R1539 VSS.n4416 VSS.n4415 292.5
R1540 VSS.n4692 VSS.n1217 292.5
R1541 VSS.n1217 VSS.n1216 292.5
R1542 VSS.n4694 VSS.n4693 292.5
R1543 VSS.n4695 VSS.n4694 292.5
R1544 VSS.n1218 VSS.n1214 292.5
R1545 VSS.n4696 VSS.n1214 292.5
R1546 VSS.n4698 VSS.n1215 292.5
R1547 VSS.n4698 VSS.n4697 292.5
R1548 VSS.n4699 VSS.n1213 292.5
R1549 VSS.n4699 VSS.n1178 292.5
R1550 VSS.n4701 VSS.n4700 292.5
R1551 VSS.n4700 VSS.n1177 292.5
R1552 VSS.n4702 VSS.n1212 292.5
R1553 VSS.n1212 VSS.n1211 292.5
R1554 VSS.n4704 VSS.n4703 292.5
R1555 VSS.n4704 VSS.n1210 292.5
R1556 VSS.n4705 VSS.n1206 292.5
R1557 VSS.n4706 VSS.n4705 292.5
R1558 VSS.n4691 VSS.n4690 292.5
R1559 VSS.n4690 VSS.n1179 292.5
R1560 VSS.n1236 VSS.n1234 292.5
R1561 VSS.n1239 VSS.n1238 292.5
R1562 VSS.n1241 VSS.n1240 292.5
R1563 VSS.n1243 VSS.n1232 292.5
R1564 VSS.n1245 VSS.n1231 292.5
R1565 VSS.n1248 VSS.n1247 292.5
R1566 VSS.n1250 VSS.n1249 292.5
R1567 VSS.n1252 VSS.n1229 292.5
R1568 VSS.n1254 VSS.n1225 292.5
R1569 VSS.n1257 VSS.n1256 292.5
R1570 VSS.n1258 VSS.n1220 292.5
R1571 VSS.n1301 VSS.n1300 292.5
R1572 VSS.n1298 VSS.n1297 292.5
R1573 VSS.n1295 VSS.n1294 292.5
R1574 VSS.n1293 VSS.n1292 292.5
R1575 VSS.n1290 VSS.n1289 292.5
R1576 VSS.n1288 VSS.n1287 292.5
R1577 VSS.n1285 VSS.n1284 292.5
R1578 VSS.n1283 VSS.n1282 292.5
R1579 VSS.n1280 VSS.n1279 292.5
R1580 VSS.n1302 VSS.n1192 292.5
R1581 VSS.n1316 VSS.n1314 292.5
R1582 VSS.n1318 VSS.n1313 292.5
R1583 VSS.n1321 VSS.n1320 292.5
R1584 VSS.n1323 VSS.n1322 292.5
R1585 VSS.n1325 VSS.n1311 292.5
R1586 VSS.n1327 VSS.n1310 292.5
R1587 VSS.n1330 VSS.n1329 292.5
R1588 VSS.n1332 VSS.n1331 292.5
R1589 VSS.n1334 VSS.n1308 292.5
R1590 VSS.n1336 VSS.n1278 292.5
R1591 VSS.n1339 VSS.n1338 292.5
R1592 VSS.n5014 VSS.n331 292.5
R1593 VSS.n5032 VSS.n5031 292.5
R1594 VSS.n5030 VSS.n5029 292.5
R1595 VSS.n5028 VSS.n5027 292.5
R1596 VSS.n5026 VSS.n5025 292.5
R1597 VSS.n5024 VSS.n5023 292.5
R1598 VSS.n5035 VSS.n5020 292.5
R1599 VSS.n5038 VSS.n5037 292.5
R1600 VSS.n5040 VSS.n5039 292.5
R1601 VSS.n5042 VSS.n5041 292.5
R1602 VSS.n4045 VSS.n4044 292.5
R1603 VSS.n4043 VSS.n4020 292.5
R1604 VSS.n4042 VSS.n4041 292.5
R1605 VSS.n4023 VSS.n4022 292.5
R1606 VSS.n4031 VSS.n4030 292.5
R1607 VSS.n4033 VSS.n4032 292.5
R1608 VSS.n4035 VSS.n4034 292.5
R1609 VSS.n4037 VSS.n4036 292.5
R1610 VSS.n4029 VSS.n4026 292.5
R1611 VSS.n4028 VSS.n4027 292.5
R1612 VSS.n4048 VSS.n4015 292.5
R1613 VSS.n3918 VSS.n3917 292.5
R1614 VSS.n3917 VSS.n1176 292.5
R1615 VSS.n3916 VSS.n3905 292.5
R1616 VSS.n3916 VSS.n3915 292.5
R1617 VSS.n3910 VSS.n3906 292.5
R1618 VSS.n3914 VSS.n3906 292.5
R1619 VSS.n3912 VSS.n3911 292.5
R1620 VSS.n3913 VSS.n3912 292.5
R1621 VSS.n3909 VSS.n3908 292.5
R1622 VSS.n3908 VSS.n3907 292.5
R1623 VSS.n1170 VSS.n1169 292.5
R1624 VSS.n1175 VSS.n1170 292.5
R1625 VSS.n4722 VSS.n4721 292.5
R1626 VSS.n4721 VSS.n4720 292.5
R1627 VSS.n4723 VSS.n1168 292.5
R1628 VSS.n1171 VSS.n1168 292.5
R1629 VSS.n4725 VSS.n4724 292.5
R1630 VSS.n4725 VSS.n1167 292.5
R1631 VSS.n4726 VSS.n1161 292.5
R1632 VSS.n4727 VSS.n4726 292.5
R1633 VSS.n3881 VSS.n3880 292.5
R1634 VSS.n3883 VSS.n3882 292.5
R1635 VSS.n3885 VSS.n3877 292.5
R1636 VSS.n3887 VSS.n3876 292.5
R1637 VSS.n3890 VSS.n3889 292.5
R1638 VSS.n3892 VSS.n3891 292.5
R1639 VSS.n3894 VSS.n3874 292.5
R1640 VSS.n3896 VSS.n3873 292.5
R1641 VSS.n3899 VSS.n3898 292.5
R1642 VSS.n3901 VSS.n3900 292.5
R1643 VSS.n3903 VSS.n3869 292.5
R1644 VSS.n3384 VSS.n3383 292.5
R1645 VSS.n3387 VSS.n3386 292.5
R1646 VSS.n3296 VSS.n3295 292.5
R1647 VSS.n3293 VSS.n3292 292.5
R1648 VSS.n3401 VSS.n3400 292.5
R1649 VSS.n3404 VSS.n3403 292.5
R1650 VSS.n3285 VSS.n3284 292.5
R1651 VSS.n3282 VSS.n3281 292.5
R1652 VSS.n3930 VSS.n3929 292.5
R1653 VSS.n3927 VSS.n3926 292.5
R1654 VSS.n3865 VSS.n3864 292.5
R1655 VSS.n3862 VSS.n3861 292.5
R1656 VSS.n3856 VSS.n3855 292.5
R1657 VSS.n3853 VSS.n3852 292.5
R1658 VSS.n3847 VSS.n3846 292.5
R1659 VSS.n3844 VSS.n3843 292.5
R1660 VSS.n1345 VSS.n1065 292.5
R1661 VSS.n1343 VSS.n1064 292.5
R1662 VSS.n4788 VSS.n4787 292.5
R1663 VSS.n4791 VSS.n4790 292.5
R1664 VSS.n2987 VSS.n2986 292.5
R1665 VSS.n2990 VSS.n2989 292.5
R1666 VSS.n2873 VSS.n2872 292.5
R1667 VSS.n2870 VSS.n2869 292.5
R1668 VSS.n3004 VSS.n3003 292.5
R1669 VSS.n3007 VSS.n3006 292.5
R1670 VSS.n2862 VSS.n2861 292.5
R1671 VSS.n2859 VSS.n2858 292.5
R1672 VSS.n3022 VSS.n3021 292.5
R1673 VSS.n3019 VSS.n3018 292.5
R1674 VSS.n2207 VSS.n1259 292.5
R1675 VSS.n2212 VSS.n2211 292.5
R1676 VSS.n2096 VSS.n2095 292.5
R1677 VSS.n2093 VSS.n2092 292.5
R1678 VSS.n2226 VSS.n2225 292.5
R1679 VSS.n2229 VSS.n2228 292.5
R1680 VSS.n2085 VSS.n2084 292.5
R1681 VSS.n2082 VSS.n2081 292.5
R1682 VSS.n2716 VSS.n2715 292.5
R1683 VSS.n2713 VSS.n2712 292.5
R1684 VSS.n3094 VSS.n3093 292.5
R1685 VSS.n3092 VSS.n3071 292.5
R1686 VSS.n3091 VSS.n3090 292.5
R1687 VSS.n3086 VSS.n3073 292.5
R1688 VSS.n3085 VSS.n3084 292.5
R1689 VSS.n3083 VSS.n3082 292.5
R1690 VSS.n3081 VSS.n3080 292.5
R1691 VSS.n3079 VSS.n3078 292.5
R1692 VSS.n3077 VSS.n3076 292.5
R1693 VSS.n3179 VSS.n1162 292.5
R1694 VSS.n3173 VSS.n3157 292.5
R1695 VSS.n3175 VSS.n3174 292.5
R1696 VSS.n3172 VSS.n3171 292.5
R1697 VSS.n3170 VSS.n3169 292.5
R1698 VSS.n3168 VSS.n3167 292.5
R1699 VSS.n3166 VSS.n3165 292.5
R1700 VSS.n3164 VSS.n3163 292.5
R1701 VSS.n3162 VSS.n3161 292.5
R1702 VSS.n3997 VSS.n3996 292.5
R1703 VSS.n3995 VSS.n3994 292.5
R1704 VSS.n3975 VSS.n3974 292.5
R1705 VSS.n3990 VSS.n3989 292.5
R1706 VSS.n3988 VSS.n3978 292.5
R1707 VSS.n3987 VSS.n3986 292.5
R1708 VSS.n3985 VSS.n3984 292.5
R1709 VSS.n3983 VSS.n3982 292.5
R1710 VSS.n3981 VSS.n3980 292.5
R1711 VSS.n4052 VSS.n4008 292.5
R1712 VSS.n4008 VSS.n1174 292.5
R1713 VSS.n4054 VSS.n4053 292.5
R1714 VSS.n4055 VSS.n4054 292.5
R1715 VSS.n4006 VSS.n4005 292.5
R1716 VSS.n4056 VSS.n4006 292.5
R1717 VSS.n4059 VSS.n4058 292.5
R1718 VSS.n4058 VSS.n4057 292.5
R1719 VSS.n4060 VSS.n4004 292.5
R1720 VSS.n4007 VSS.n4004 292.5
R1721 VSS.n4062 VSS.n4061 292.5
R1722 VSS.n4062 VSS.n1173 292.5
R1723 VSS.n4063 VSS.n4003 292.5
R1724 VSS.n4063 VSS.n1172 292.5
R1725 VSS.n4066 VSS.n4065 292.5
R1726 VSS.n4065 VSS.n4064 292.5
R1727 VSS.n4067 VSS.n4002 292.5
R1728 VSS.n4002 VSS.n4001 292.5
R1729 VSS.n4069 VSS.n4068 292.5
R1730 VSS.n4070 VSS.n4069 292.5
R1731 VSS.n2769 VSS.n1207 292.5
R1732 VSS.n2769 VSS.n2768 292.5
R1733 VSS.n2772 VSS.n2770 292.5
R1734 VSS.n2770 VSS.n2766 292.5
R1735 VSS.n2774 VSS.n2773 292.5
R1736 VSS.n2775 VSS.n2774 292.5
R1737 VSS.n2771 VSS.n2764 292.5
R1738 VSS.n2776 VSS.n2764 292.5
R1739 VSS.n2778 VSS.n2765 292.5
R1740 VSS.n2778 VSS.n2777 292.5
R1741 VSS.n2779 VSS.n2763 292.5
R1742 VSS.n2780 VSS.n2779 292.5
R1743 VSS.n2783 VSS.n2782 292.5
R1744 VSS.n2782 VSS.n2781 292.5
R1745 VSS.n2784 VSS.n2762 292.5
R1746 VSS.n2762 VSS.n2761 292.5
R1747 VSS.n2786 VSS.n2785 292.5
R1748 VSS.n2787 VSS.n2786 292.5
R1749 VSS.n2788 VSS.n2037 292.5
R1750 VSS.n2790 VSS.n2789 292.5
R1751 VSS.n2767 VSS.n1205 292.5
R1752 VSS.n4214 VSS.n4213 292.5
R1753 VSS.n4217 VSS.n4216 292.5
R1754 VSS.n4223 VSS.n4222 292.5
R1755 VSS.n4226 VSS.n4225 292.5
R1756 VSS.n4235 VSS.n4234 292.5
R1757 VSS.n4238 VSS.n4237 292.5
R1758 VSS.n4247 VSS.n4246 292.5
R1759 VSS.n4249 VSS.n1840 292.5
R1760 VSS.n4251 VSS.n1811 292.5
R1761 VSS.n4253 VSS.n1810 292.5
R1762 VSS.n4256 VSS.n4255 292.5
R1763 VSS.n1836 VSS.n1833 292.5
R1764 VSS.n3971 VSS.n3970 292.5
R1765 VSS.n3968 VSS.n3967 292.5
R1766 VSS.n3339 VSS.n3338 292.5
R1767 VSS.n3336 VSS.n3307 292.5
R1768 VSS.n3334 VSS.n3333 292.5
R1769 VSS.n3311 VSS.n3310 292.5
R1770 VSS.n3313 VSS.n3309 292.5
R1771 VSS.n3316 VSS.n3315 292.5
R1772 VSS.n3957 VSS.n3956 292.5
R1773 VSS.n3960 VSS.n3959 292.5
R1774 VSS.n3270 VSS.n3269 292.5
R1775 VSS.n3267 VSS.n1164 292.5
R1776 VSS.n4734 VSS.n4733 292.5
R1777 VSS.n4737 VSS.n4736 292.5
R1778 VSS.n1156 VSS.n1151 292.5
R1779 VSS.n1154 VSS.n1150 292.5
R1780 VSS.n4747 VSS.n4746 292.5
R1781 VSS.n4750 VSS.n4749 292.5
R1782 VSS.n1140 VSS.n1136 292.5
R1783 VSS.n1138 VSS.n1135 292.5
R1784 VSS.n4760 VSS.n4759 292.5
R1785 VSS.n4762 VSS.n1089 292.5
R1786 VSS.n4764 VSS.n1088 292.5
R1787 VSS.n4767 VSS.n4766 292.5
R1788 VSS.n1197 VSS.n1194 292.5
R1789 VSS.n2939 VSS.n2938 292.5
R1790 VSS.n2935 VSS.n2904 292.5
R1791 VSS.n2933 VSS.n2903 292.5
R1792 VSS.n2931 VSS.n2930 292.5
R1793 VSS.n2908 VSS.n2907 292.5
R1794 VSS.n2910 VSS.n2906 292.5
R1795 VSS.n2913 VSS.n2912 292.5
R1796 VSS.n3049 VSS.n3048 292.5
R1797 VSS.n3052 VSS.n3051 292.5
R1798 VSS.n2847 VSS.n2846 292.5
R1799 VSS.n2844 VSS.n1209 292.5
R1800 VSS.n1203 VSS.n1201 292.5
R1801 VSS.n2160 VSS.n2159 292.5
R1802 VSS.n2156 VSS.n2125 292.5
R1803 VSS.n2154 VSS.n2124 292.5
R1804 VSS.n2152 VSS.n2151 292.5
R1805 VSS.n2129 VSS.n2128 292.5
R1806 VSS.n2131 VSS.n2127 292.5
R1807 VSS.n2134 VSS.n2133 292.5
R1808 VSS.n2743 VSS.n2742 292.5
R1809 VSS.n2746 VSS.n2745 292.5
R1810 VSS.n2679 VSS.n2678 292.5
R1811 VSS.n2682 VSS.n2681 292.5
R1812 VSS.n4707 VSS.n1208 292.5
R1813 VSS.n4728 VSS.n1163 292.5
R1814 VSS.n4071 VSS.n3999 292.5
R1815 VSS.n2489 VSS.n1356 292.5
R1816 VSS.n2484 VSS.n2483 292.5
R1817 VSS.n2478 VSS.n2477 292.5
R1818 VSS.n2475 VSS.n2474 292.5
R1819 VSS.n2469 VSS.n2468 292.5
R1820 VSS.n2466 VSS.n2465 292.5
R1821 VSS.n1789 VSS.n1788 292.5
R1822 VSS.n1786 VSS.n1785 292.5
R1823 VSS.n4292 VSS.n4291 292.5
R1824 VSS.n4295 VSS.n4294 292.5
R1825 VSS.n2515 VSS.n2514 292.5
R1826 VSS.n2512 VSS.n2511 292.5
R1827 VSS.n2414 VSS.n2411 292.5
R1828 VSS.n2416 VSS.n2412 292.5
R1829 VSS.n2418 VSS.n2413 292.5
R1830 VSS.n2421 VSS.n2420 292.5
R1831 VSS.n4349 VSS.n4348 292.5
R1832 VSS.n4351 VSS.n1759 292.5
R1833 VSS.n4354 VSS.n4353 292.5
R1834 VSS.n4315 VSS.n1752 292.5
R1835 VSS.n4317 VSS.n1751 292.5
R1836 VSS.n4320 VSS.n4319 292.5
R1837 VSS.n4422 VSS.n4421 292.5
R1838 VSS.n4425 VSS.n4424 292.5
R1839 VSS.n1559 VSS.n1554 292.5
R1840 VSS.n1557 VSS.n1553 292.5
R1841 VSS.n4435 VSS.n4434 292.5
R1842 VSS.n4438 VSS.n4437 292.5
R1843 VSS.n1543 VSS.n1539 292.5
R1844 VSS.n1541 VSS.n1538 292.5
R1845 VSS.n4448 VSS.n4447 292.5
R1846 VSS.n4450 VSS.n1511 292.5
R1847 VSS.n4452 VSS.n1510 292.5
R1848 VSS.n4455 VSS.n4454 292.5
R1849 VSS.n737 VSS.n735 292.5
R1850 VSS.n3810 VSS.n3809 292.5
R1851 VSS.n3806 VSS.n3805 292.5
R1852 VSS.n3766 VSS.n3756 292.5
R1853 VSS.n3768 VSS.n3757 292.5
R1854 VSS.n3770 VSS.n3765 292.5
R1855 VSS.n3772 VSS.n3758 292.5
R1856 VSS.n3774 VSS.n3759 292.5
R1857 VSS.n3777 VSS.n3776 292.5
R1858 VSS.n3763 VSS.n1032 292.5
R1859 VSS.n3761 VSS.n1031 292.5
R1860 VSS.n731 VSS.n730 292.5
R1861 VSS.n5048 VSS.n5047 292.5
R1862 VSS.n5051 VSS.n5050 292.5
R1863 VSS.n722 VSS.n717 292.5
R1864 VSS.n720 VSS.n716 292.5
R1865 VSS.n5061 VSS.n5060 292.5
R1866 VSS.n5064 VSS.n5063 292.5
R1867 VSS.n706 VSS.n702 292.5
R1868 VSS.n704 VSS.n701 292.5
R1869 VSS.n5074 VSS.n5073 292.5
R1870 VSS.n5076 VSS.n491 292.5
R1871 VSS.n5078 VSS.n490 292.5
R1872 VSS.n5081 VSS.n5080 292.5
R1873 VSS.n5255 VSS.n5254 292.5
R1874 VSS.n5258 VSS.n5257 292.5
R1875 VSS.n294 VSS.n289 292.5
R1876 VSS.n292 VSS.n288 292.5
R1877 VSS.n5268 VSS.n5267 292.5
R1878 VSS.n5271 VSS.n5270 292.5
R1879 VSS.n278 VSS.n274 292.5
R1880 VSS.n276 VSS.n273 292.5
R1881 VSS.n5281 VSS.n5280 292.5
R1882 VSS.n5283 VSS.n242 292.5
R1883 VSS.n5285 VSS.n241 292.5
R1884 VSS.n5288 VSS.n5287 292.5
R1885 VSS.n5466 VSS.n5465 292.5
R1886 VSS.n5460 VSS.n63 292.5
R1887 VSS.n5459 VSS.n5458 292.5
R1888 VSS.n5457 VSS.n5456 292.5
R1889 VSS.n5455 VSS.n5454 292.5
R1890 VSS.n5452 VSS.n5451 292.5
R1891 VSS.n5450 VSS.n5449 292.5
R1892 VSS.n5447 VSS.n5446 292.5
R1893 VSS.n5445 VSS.n5444 292.5
R1894 VSS.n5442 VSS.n5441 292.5
R1895 VSS.n5440 VSS.n5439 292.5
R1896 VSS.n4618 VSS.n1373 292.5
R1897 VSS.t79 VSS.n4618 292.5
R1898 VSS.n4619 VSS.n1372 292.5
R1899 VSS.n4619 VSS.t79 292.5
R1900 VSS.n4677 VSS.n1265 284.909
R1901 VSS.n4641 VSS.n4640 284.909
R1902 VSS.n5539 VSS.n20 284.909
R1903 VSS.n1887 VSS.t75 284.663
R1904 VSS.n1882 VSS.t62 284.339
R1905 VSS.n5222 VSS.n358 272.089
R1906 VSS.n5224 VSS.n341 272.089
R1907 VSS.n358 VSS.n357 272.089
R1908 VSS.n5224 VSS.n340 272.089
R1909 VSS.n358 VSS.n345 272.089
R1910 VSS.n5224 VSS.n339 272.089
R1911 VSS.n358 VSS.n344 272.089
R1912 VSS.n5225 VSS.n5224 272.089
R1913 VSS.n358 VSS.n336 272.089
R1914 VSS.n5224 VSS.n338 272.089
R1915 VSS.n5215 VSS.n366 272.089
R1916 VSS.n389 VSS.n388 272.089
R1917 VSS.n5215 VSS.n365 272.089
R1918 VSS.n388 VSS.n387 272.089
R1919 VSS.n5215 VSS.n364 272.089
R1920 VSS.n388 VSS.n372 272.089
R1921 VSS.n5215 VSS.n363 272.089
R1922 VSS.n388 VSS.n371 272.089
R1923 VSS.n5215 VSS.n362 272.089
R1924 VSS.n388 VSS.n360 272.089
R1925 VSS.n4962 VSS.n781 272.089
R1926 VSS.n804 VSS.n803 272.089
R1927 VSS.n4962 VSS.n780 272.089
R1928 VSS.n803 VSS.n802 272.089
R1929 VSS.n4962 VSS.n779 272.089
R1930 VSS.n803 VSS.n787 272.089
R1931 VSS.n4962 VSS.n778 272.089
R1932 VSS.n803 VSS.n786 272.089
R1933 VSS.n4962 VSS.n777 272.089
R1934 VSS.n803 VSS.n775 272.089
R1935 VSS.n2360 VSS.n209 272.089
R1936 VSS.n5322 VSS.n209 272.089
R1937 VSS.n212 VSS.n209 272.089
R1938 VSS.n620 VSS.n209 272.089
R1939 VSS.n634 VSS.n209 272.089
R1940 VSS.n642 VSS.n209 272.089
R1941 VSS.n465 VSS.n209 272.089
R1942 VSS.n466 VSS.n209 272.089
R1943 VSS.n916 VSS.n209 272.089
R1944 VSS.n912 VSS.n209 272.089
R1945 VSS.n938 VSS.n209 272.089
R1946 VSS.n333 VSS.n209 272.089
R1947 VSS.n1006 VSS.n209 272.089
R1948 VSS.n1007 VSS.n209 272.089
R1949 VSS.n3711 VSS.n209 272.089
R1950 VSS.n3707 VSS.n209 272.089
R1951 VSS.n3733 VSS.n209 272.089
R1952 VSS.n762 VSS.n209 272.089
R1953 VSS.n1485 VSS.n209 272.089
R1954 VSS.n1486 VSS.n209 272.089
R1955 VSS.n1625 VSS.n209 272.089
R1956 VSS.n1621 VSS.n209 272.089
R1957 VSS.n1647 VSS.n209 272.089
R1958 VSS.n1688 VSS.n209 272.089
R1959 VSS.n4373 VSS.n209 272.089
R1960 VSS.n1700 VSS.n209 272.089
R1961 VSS.n1712 VSS.n209 272.089
R1962 VSS.n1733 VSS.n209 272.089
R1963 VSS.n1731 VSS.n211 272.089
R1964 VSS.n1730 VSS.n211 272.089
R1965 VSS.n1715 VSS.n211 272.089
R1966 VSS.n4371 VSS.n211 272.089
R1967 VSS.n1698 VSS.n211 272.089
R1968 VSS.n4400 VSS.n211 272.089
R1969 VSS.n1646 VSS.n211 272.089
R1970 VSS.n1637 VSS.n211 272.089
R1971 VSS.n1628 VSS.n211 272.089
R1972 VSS.n4487 VSS.n211 272.089
R1973 VSS.n1483 VSS.n211 272.089
R1974 VSS.n3732 VSS.n211 272.089
R1975 VSS.n3723 VSS.n211 272.089
R1976 VSS.n3714 VSS.n211 272.089
R1977 VSS.n4860 VSS.n211 272.089
R1978 VSS.n1004 VSS.n211 272.089
R1979 VSS.n937 VSS.n211 272.089
R1980 VSS.n928 VSS.n211 272.089
R1981 VSS.n919 VSS.n211 272.089
R1982 VSS.n5113 VSS.n211 272.089
R1983 VSS.n640 VSS.n211 272.089
R1984 VSS.n635 VSS.n211 272.089
R1985 VSS.n615 VSS.n211 272.089
R1986 VSS.n618 VSS.n211 272.089
R1987 VSS.n5320 VSS.n211 272.089
R1988 VSS.n211 VSS.n208 272.089
R1989 VSS.n2362 VSS.n211 272.089
R1990 VSS.n2281 VSS.n23 272.089
R1991 VSS.n5342 VSS.n23 272.089
R1992 VSS.n179 VSS.n23 272.089
R1993 VSS.n582 VSS.n23 272.089
R1994 VSS.n591 VSS.n23 272.089
R1995 VSS.n84 VSS.n23 272.089
R1996 VSS.n434 VSS.n23 272.089
R1997 VSS.n435 VSS.n23 272.089
R1998 VSS.n855 VSS.n23 272.089
R1999 VSS.n870 VSS.n23 272.089
R2000 VSS.n964 VSS.n23 272.089
R2001 VSS.n968 VSS.n23 272.089
R2002 VSS.n972 VSS.n23 272.089
R2003 VSS.n973 VSS.n23 272.089
R2004 VSS.n3455 VSS.n23 272.089
R2005 VSS.n3451 VSS.n23 272.089
R2006 VSS.n3682 VSS.n23 272.089
R2007 VSS.n3678 VSS.n23 272.089
R2008 VSS.n3480 VSS.n23 272.089
R2009 VSS.n3519 VSS.n23 272.089
R2010 VSS.n3553 VSS.n23 272.089
R2011 VSS.n3535 VSS.n23 272.089
R2012 VSS.n3541 VSS.n23 272.089
R2013 VSS.n1446 VSS.n23 272.089
R2014 VSS.n1447 VSS.n23 272.089
R2015 VSS.n4561 VSS.n23 272.089
R2016 VSS.n4534 VSS.n23 272.089
R2017 VSS.n26 VSS.n23 272.089
R2018 VSS.n5534 VSS.n25 272.089
R2019 VSS.n4546 VSS.n25 272.089
R2020 VSS.n4559 VSS.n25 272.089
R2021 VSS.n4532 VSS.n25 272.089
R2022 VSS.n4574 VSS.n25 272.089
R2023 VSS.n4503 VSS.n25 272.089
R2024 VSS.n3543 VSS.n25 272.089
R2025 VSS.n3551 VSS.n25 272.089
R2026 VSS.n3534 VSS.n25 272.089
R2027 VSS.n3525 VSS.n25 272.089
R2028 VSS.n3676 VSS.n25 272.089
R2029 VSS.n3475 VSS.n25 272.089
R2030 VSS.n3466 VSS.n25 272.089
R2031 VSS.n3457 VSS.n25 272.089
R2032 VSS.n4879 VSS.n25 272.089
R2033 VSS.n970 VSS.n25 272.089
R2034 VSS.n848 VSS.n25 272.089
R2035 VSS.n850 VSS.n25 272.089
R2036 VSS.n853 VSS.n25 272.089
R2037 VSS.n5132 VSS.n25 272.089
R2038 VSS.n432 VSS.n25 272.089
R2039 VSS.n592 VSS.n25 272.089
R2040 VSS.n569 VSS.n25 272.089
R2041 VSS.n572 VSS.n25 272.089
R2042 VSS.n5340 VSS.n25 272.089
R2043 VSS.n177 VSS.n25 272.089
R2044 VSS.n2283 VSS.n25 272.089
R2045 VSS.n5428 VSS.n92 272.089
R2046 VSS.n157 VSS.n156 272.089
R2047 VSS.n5428 VSS.n91 272.089
R2048 VSS.n157 VSS.n137 272.089
R2049 VSS.n5428 VSS.n90 272.089
R2050 VSS.n157 VSS.n136 272.089
R2051 VSS.n5428 VSS.n89 272.089
R2052 VSS.n157 VSS.n135 272.089
R2053 VSS.n5428 VSS.n88 272.089
R2054 VSS.n157 VSS.n86 272.089
R2055 VSS.n5241 VSS.n5240 272.089
R2056 VSS.n5251 VSS.n304 272.089
R2057 VSS.n5241 VSS.n311 272.089
R2058 VSS.n5251 VSS.n305 272.089
R2059 VSS.n5241 VSS.n310 272.089
R2060 VSS.n5251 VSS.n306 272.089
R2061 VSS.n5243 VSS.n5241 272.089
R2062 VSS.n5251 VSS.n307 272.089
R2063 VSS.n5241 VSS.n308 272.089
R2064 VSS.n5251 VSS.n5250 272.089
R2065 VSS.n4997 VSS.n4996 272.089
R2066 VSS.n5007 VSS.n744 272.089
R2067 VSS.n4997 VSS.n751 272.089
R2068 VSS.n5007 VSS.n745 272.089
R2069 VSS.n4997 VSS.n750 272.089
R2070 VSS.n5007 VSS.n746 272.089
R2071 VSS.n4999 VSS.n4997 272.089
R2072 VSS.n5007 VSS.n747 272.089
R2073 VSS.n4997 VSS.n748 272.089
R2074 VSS.n5007 VSS.n5006 272.089
R2075 VSS.n4408 VSS.n4407 272.089
R2076 VSS.n4418 VSS.n1568 272.089
R2077 VSS.n4408 VSS.n1575 272.089
R2078 VSS.n4418 VSS.n1569 272.089
R2079 VSS.n4408 VSS.n1574 272.089
R2080 VSS.n4418 VSS.n1570 272.089
R2081 VSS.n4410 VSS.n4408 272.089
R2082 VSS.n4418 VSS.n1571 272.089
R2083 VSS.n4408 VSS.n1572 272.089
R2084 VSS.n4418 VSS.n4417 272.089
R2085 VSS.n1235 VSS.n1228 272.089
R2086 VSS.n1237 VSS.n1227 272.089
R2087 VSS.n1233 VSS.n1228 272.089
R2088 VSS.n1242 VSS.n1227 272.089
R2089 VSS.n1244 VSS.n1228 272.089
R2090 VSS.n1246 VSS.n1227 272.089
R2091 VSS.n1230 VSS.n1228 272.089
R2092 VSS.n1251 VSS.n1227 272.089
R2093 VSS.n1253 VSS.n1228 272.089
R2094 VSS.n1255 VSS.n1227 272.089
R2095 VSS.n1228 VSS.n1226 272.089
R2096 VSS.n4719 VSS.n1191 272.089
R2097 VSS.n1296 VSS.n1186 272.089
R2098 VSS.n4719 VSS.n1190 272.089
R2099 VSS.n1291 VSS.n1186 272.089
R2100 VSS.n4719 VSS.n1189 272.089
R2101 VSS.n1286 VSS.n1186 272.089
R2102 VSS.n4719 VSS.n1188 272.089
R2103 VSS.n1281 VSS.n1186 272.089
R2104 VSS.n4719 VSS.n1187 272.089
R2105 VSS.n1299 VSS.n1186 272.089
R2106 VSS.n1317 VSS.n1306 272.089
R2107 VSS.n1315 VSS.n1307 272.089
R2108 VSS.n1319 VSS.n1307 272.089
R2109 VSS.n1312 VSS.n1306 272.089
R2110 VSS.n1324 VSS.n1307 272.089
R2111 VSS.n1326 VSS.n1306 272.089
R2112 VSS.n1328 VSS.n1307 272.089
R2113 VSS.n1309 VSS.n1306 272.089
R2114 VSS.n1333 VSS.n1307 272.089
R2115 VSS.n1335 VSS.n1306 272.089
R2116 VSS.n1337 VSS.n1307 272.089
R2117 VSS.n5034 VSS.n5033 272.089
R2118 VSS.n5044 VSS.n5015 272.089
R2119 VSS.n5034 VSS.n5022 272.089
R2120 VSS.n5044 VSS.n5016 272.089
R2121 VSS.n5034 VSS.n5021 272.089
R2122 VSS.n5044 VSS.n5017 272.089
R2123 VSS.n5036 VSS.n5034 272.089
R2124 VSS.n5044 VSS.n5018 272.089
R2125 VSS.n5034 VSS.n5019 272.089
R2126 VSS.n5044 VSS.n5043 272.089
R2127 VSS.n4039 VSS.n4021 272.089
R2128 VSS.n4047 VSS.n4046 272.089
R2129 VSS.n4040 VSS.n4039 272.089
R2130 VSS.n4047 VSS.n4019 272.089
R2131 VSS.n4039 VSS.n4024 272.089
R2132 VSS.n4047 VSS.n4018 272.089
R2133 VSS.n4039 VSS.n4025 272.089
R2134 VSS.n4047 VSS.n4017 272.089
R2135 VSS.n4039 VSS.n4038 272.089
R2136 VSS.n4047 VSS.n4016 272.089
R2137 VSS.n4039 VSS.n4012 272.089
R2138 VSS.n3878 VSS.n3870 272.089
R2139 VSS.n3879 VSS.n3871 272.089
R2140 VSS.n3884 VSS.n3871 272.089
R2141 VSS.n3886 VSS.n3870 272.089
R2142 VSS.n3888 VSS.n3871 272.089
R2143 VSS.n3875 VSS.n3870 272.089
R2144 VSS.n3893 VSS.n3871 272.089
R2145 VSS.n3895 VSS.n3870 272.089
R2146 VSS.n3897 VSS.n3871 272.089
R2147 VSS.n3872 VSS.n3870 272.089
R2148 VSS.n3902 VSS.n3871 272.089
R2149 VSS.n4683 VSS.n1266 272.089
R2150 VSS.n4683 VSS.n1267 272.089
R2151 VSS.n4683 VSS.n1268 272.089
R2152 VSS.n4683 VSS.n1269 272.089
R2153 VSS.n4683 VSS.n1270 272.089
R2154 VSS.n4684 VSS.n4683 272.089
R2155 VSS.n4683 VSS.n1222 272.089
R2156 VSS.n4683 VSS.n1271 272.089
R2157 VSS.n4683 VSS.n1272 272.089
R2158 VSS.n4683 VSS.n1273 272.089
R2159 VSS.n4683 VSS.n1274 272.089
R2160 VSS.n4683 VSS.n1342 272.089
R2161 VSS.n4683 VSS.n1059 272.089
R2162 VSS.n4683 VSS.n1061 272.089
R2163 VSS.n4683 VSS.n1346 272.089
R2164 VSS.n4683 VSS.n1347 272.089
R2165 VSS.n4683 VSS.n1348 272.089
R2166 VSS.n4683 VSS.n1349 272.089
R2167 VSS.n4683 VSS.n1350 272.089
R2168 VSS.n4683 VSS.n1351 272.089
R2169 VSS.n4683 VSS.n1352 272.089
R2170 VSS.n4683 VSS.n1353 272.089
R2171 VSS.n4683 VSS.n1354 272.089
R2172 VSS.n4683 VSS.n1355 272.089
R2173 VSS.n4683 VSS.n4682 272.089
R2174 VSS.n3385 VSS.n1060 272.089
R2175 VSS.n3294 VSS.n1060 272.089
R2176 VSS.n3402 VSS.n1060 272.089
R2177 VSS.n3283 VSS.n1060 272.089
R2178 VSS.n3928 VSS.n1060 272.089
R2179 VSS.n3863 VSS.n1060 272.089
R2180 VSS.n3854 VSS.n1060 272.089
R2181 VSS.n3845 VSS.n1060 272.089
R2182 VSS.n1344 VSS.n1060 272.089
R2183 VSS.n4789 VSS.n1060 272.089
R2184 VSS.n2988 VSS.n1060 272.089
R2185 VSS.n2871 VSS.n1060 272.089
R2186 VSS.n3005 VSS.n1060 272.089
R2187 VSS.n2860 VSS.n1060 272.089
R2188 VSS.n3020 VSS.n1060 272.089
R2189 VSS.n2210 VSS.n1060 272.089
R2190 VSS.n2094 VSS.n1060 272.089
R2191 VSS.n2227 VSS.n1060 272.089
R2192 VSS.n2083 VSS.n1060 272.089
R2193 VSS.n2714 VSS.n1060 272.089
R2194 VSS.n3096 VSS.n3095 272.089
R2195 VSS.n3089 VSS.n3088 272.089
R2196 VSS.n3096 VSS.n3070 272.089
R2197 VSS.n3088 VSS.n3087 272.089
R2198 VSS.n3096 VSS.n3069 272.089
R2199 VSS.n3088 VSS.n3075 272.089
R2200 VSS.n3096 VSS.n3068 272.089
R2201 VSS.n3088 VSS.n3074 272.089
R2202 VSS.n3096 VSS.n3067 272.089
R2203 VSS.n3181 VSS.n3180 272.089
R2204 VSS.n3177 VSS.n3176 272.089
R2205 VSS.n3181 VSS.n3156 272.089
R2206 VSS.n3177 VSS.n3160 272.089
R2207 VSS.n3181 VSS.n3155 272.089
R2208 VSS.n3177 VSS.n3159 272.089
R2209 VSS.n3181 VSS.n3154 272.089
R2210 VSS.n3177 VSS.n3158 272.089
R2211 VSS.n3181 VSS.n3153 272.089
R2212 VSS.n4075 VSS.n1920 272.089
R2213 VSS.n3993 VSS.n3992 272.089
R2214 VSS.n4075 VSS.n1919 272.089
R2215 VSS.n3992 VSS.n3991 272.089
R2216 VSS.n4075 VSS.n1918 272.089
R2217 VSS.n3992 VSS.n3977 272.089
R2218 VSS.n4075 VSS.n1917 272.089
R2219 VSS.n3992 VSS.n3976 272.089
R2220 VSS.n4075 VSS.n1916 272.089
R2221 VSS.n2760 VSS.n2759 272.089
R2222 VSS.n3088 VSS.n3066 272.089
R2223 VSS.n3177 VSS.n3152 272.089
R2224 VSS.n3992 VSS.n1914 272.089
R2225 VSS.n3088 VSS.n3072 272.089
R2226 VSS.n3178 VSS.n3177 272.089
R2227 VSS.n3992 VSS.n1921 272.089
R2228 VSS.n2066 VSS.n1131 272.089
R2229 VSS.n2067 VSS.n1131 272.089
R2230 VSS.n2130 VSS.n1131 272.089
R2231 VSS.n2153 VSS.n1131 272.089
R2232 VSS.n2157 VSS.n1131 272.089
R2233 VSS.n2023 VSS.n1131 272.089
R2234 VSS.n2024 VSS.n1131 272.089
R2235 VSS.n2909 VSS.n1131 272.089
R2236 VSS.n2932 VSS.n1131 272.089
R2237 VSS.n2936 VSS.n1131 272.089
R2238 VSS.n4763 VSS.n1131 272.089
R2239 VSS.n1133 VSS.n1131 272.089
R2240 VSS.n1141 VSS.n1131 272.089
R2241 VSS.n1142 VSS.n1131 272.089
R2242 VSS.n1157 VSS.n1131 272.089
R2243 VSS.n1947 VSS.n1131 272.089
R2244 VSS.n1948 VSS.n1131 272.089
R2245 VSS.n3312 VSS.n1131 272.089
R2246 VSS.n3335 VSS.n1131 272.089
R2247 VSS.n1923 VSS.n1131 272.089
R2248 VSS.n4254 VSS.n1131 272.089
R2249 VSS.n4250 VSS.n1131 272.089
R2250 VSS.n1841 VSS.n1131 272.089
R2251 VSS.n1843 VSS.n1131 272.089
R2252 VSS.n1847 VSS.n1131 272.089
R2253 VSS.n4215 VSS.n1132 272.089
R2254 VSS.n4224 VSS.n1132 272.089
R2255 VSS.n4236 VSS.n1132 272.089
R2256 VSS.n4248 VSS.n1132 272.089
R2257 VSS.n4252 VSS.n1132 272.089
R2258 VSS.n1837 VSS.n1132 272.089
R2259 VSS.n3969 VSS.n1132 272.089
R2260 VSS.n3337 VSS.n1132 272.089
R2261 VSS.n3308 VSS.n1132 272.089
R2262 VSS.n3314 VSS.n1132 272.089
R2263 VSS.n3958 VSS.n1132 272.089
R2264 VSS.n3268 VSS.n1132 272.089
R2265 VSS.n4735 VSS.n1132 272.089
R2266 VSS.n1155 VSS.n1132 272.089
R2267 VSS.n4748 VSS.n1132 272.089
R2268 VSS.n1139 VSS.n1132 272.089
R2269 VSS.n4761 VSS.n1132 272.089
R2270 VSS.n4765 VSS.n1132 272.089
R2271 VSS.n2937 VSS.n1132 272.089
R2272 VSS.n2934 VSS.n1132 272.089
R2273 VSS.n2905 VSS.n1132 272.089
R2274 VSS.n2911 VSS.n1132 272.089
R2275 VSS.n3050 VSS.n1132 272.089
R2276 VSS.n2845 VSS.n1132 272.089
R2277 VSS.n2158 VSS.n1132 272.089
R2278 VSS.n2155 VSS.n1132 272.089
R2279 VSS.n2126 VSS.n1132 272.089
R2280 VSS.n2132 VSS.n1132 272.089
R2281 VSS.n2744 VSS.n1132 272.089
R2282 VSS.n2680 VSS.n1132 272.089
R2283 VSS.n4711 VSS.n1204 272.089
R2284 VSS.n4717 VSS.n1186 272.089
R2285 VSS.n4732 VSS.n1159 272.089
R2286 VSS.n4000 VSS.n3972 272.089
R2287 VSS.n4683 VSS.n1264 272.089
R2288 VSS.n4683 VSS.n1263 272.089
R2289 VSS.n4683 VSS.n1262 272.089
R2290 VSS.n4683 VSS.n1261 272.089
R2291 VSS.n4683 VSS.n1260 272.089
R2292 VSS.n2482 VSS.n1060 272.089
R2293 VSS.n2476 VSS.n1060 272.089
R2294 VSS.n2467 VSS.n1060 272.089
R2295 VSS.n1787 VSS.n1060 272.089
R2296 VSS.n4293 VSS.n1060 272.089
R2297 VSS.n5284 VSS.n269 272.089
R2298 VSS.n271 VSS.n269 272.089
R2299 VSS.n279 VSS.n269 272.089
R2300 VSS.n280 VSS.n269 272.089
R2301 VSS.n295 VSS.n269 272.089
R2302 VSS.n5077 VSS.n269 272.089
R2303 VSS.n699 VSS.n269 272.089
R2304 VSS.n707 VSS.n269 272.089
R2305 VSS.n708 VSS.n269 272.089
R2306 VSS.n723 VSS.n269 272.089
R2307 VSS.n3762 VSS.n269 272.089
R2308 VSS.n3775 VSS.n269 272.089
R2309 VSS.n3771 VSS.n269 272.089
R2310 VSS.n3767 VSS.n269 272.089
R2311 VSS.n3807 VSS.n269 272.089
R2312 VSS.n4451 VSS.n269 272.089
R2313 VSS.n1536 VSS.n269 272.089
R2314 VSS.n1544 VSS.n269 272.089
R2315 VSS.n1545 VSS.n269 272.089
R2316 VSS.n1560 VSS.n269 272.089
R2317 VSS.n4316 VSS.n269 272.089
R2318 VSS.n4352 VSS.n269 272.089
R2319 VSS.n1760 VSS.n269 272.089
R2320 VSS.n2417 VSS.n269 272.089
R2321 VSS.n2410 VSS.n269 272.089
R2322 VSS.n2513 VSS.n270 272.089
R2323 VSS.n2415 VSS.n270 272.089
R2324 VSS.n2419 VSS.n270 272.089
R2325 VSS.n4350 VSS.n270 272.089
R2326 VSS.n1758 VSS.n270 272.089
R2327 VSS.n4318 VSS.n270 272.089
R2328 VSS.n4423 VSS.n270 272.089
R2329 VSS.n1558 VSS.n270 272.089
R2330 VSS.n4436 VSS.n270 272.089
R2331 VSS.n1542 VSS.n270 272.089
R2332 VSS.n4449 VSS.n270 272.089
R2333 VSS.n4453 VSS.n270 272.089
R2334 VSS.n3808 VSS.n270 272.089
R2335 VSS.n3755 VSS.n270 272.089
R2336 VSS.n3769 VSS.n270 272.089
R2337 VSS.n3773 VSS.n270 272.089
R2338 VSS.n3764 VSS.n270 272.089
R2339 VSS.n3760 VSS.n270 272.089
R2340 VSS.n5049 VSS.n270 272.089
R2341 VSS.n721 VSS.n270 272.089
R2342 VSS.n5062 VSS.n270 272.089
R2343 VSS.n705 VSS.n270 272.089
R2344 VSS.n5075 VSS.n270 272.089
R2345 VSS.n5079 VSS.n270 272.089
R2346 VSS.n5256 VSS.n270 272.089
R2347 VSS.n293 VSS.n270 272.089
R2348 VSS.n5269 VSS.n270 272.089
R2349 VSS.n277 VSS.n270 272.089
R2350 VSS.n5282 VSS.n270 272.089
R2351 VSS.n5286 VSS.n270 272.089
R2352 VSS.n5241 VSS.n301 272.089
R2353 VSS.n5034 VSS.n729 272.089
R2354 VSS.n4997 VSS.n741 272.089
R2355 VSS.n4408 VSS.n1565 272.089
R2356 VSS.n157 VSS.n93 272.089
R2357 VSS.n388 VSS.n367 272.089
R2358 VSS.n803 VSS.n782 272.089
R2359 VSS.n5464 VSS.n5462 272.089
R2360 VSS.n64 VSS.n13 272.089
R2361 VSS.n5462 VSS.n5461 272.089
R2362 VSS.n69 VSS.n13 272.089
R2363 VSS.n5462 VSS.n68 272.089
R2364 VSS.n5453 VSS.n13 272.089
R2365 VSS.n5462 VSS.n67 272.089
R2366 VSS.n5448 VSS.n13 272.089
R2367 VSS.n5462 VSS.n66 272.089
R2368 VSS.n5443 VSS.n13 272.089
R2369 VSS.n5462 VSS.n65 272.089
R2370 VSS.n5468 VSS.n59 272.089
R2371 VSS.n4954 VSS.n783 272.089
R2372 VSS.n5207 VSS.n368 272.089
R2373 VSS.n5420 VSS.n94 272.089
R2374 VSS.n2547 VSS.n2546 270.175
R2375 VSS.n5374 VSS.n167 264.301
R2376 VSS.n2683 VSS.n2583 264.301
R2377 VSS.n2252 VSS.n267 264.301
R2378 VSS.n2365 VSS.n2264 264.301
R2379 VSS.n2300 VSS.n2299 264.301
R2380 VSS.n4212 VSS.n1852 264.301
R2381 VSS.n2520 VSS.n2516 264.301
R2382 VSS.n5561 VSS.n6 264.301
R2383 VSS.n4151 VSS.n1869 259.416
R2384 VSS.n1781 VSS.n1777 258.334
R2385 VSS.n4096 VSS.n4095 258.334
R2386 VSS.n3250 VSS.n3249 258.334
R2387 VSS.n3108 VSS.n3107 258.334
R2388 VSS.n2827 VSS.n2826 258.334
R2389 VSS.n1057 VSS.n1053 258.334
R2390 VSS.n4779 VSS.n1086 258.334
R2391 VSS.n5310 VSS.n239 258.334
R2392 VSS.n5351 VSS.n5350 258.334
R2393 VSS.n5330 VSS.n200 258.334
R2394 VSS.n5141 VSS.n5140 258.334
R2395 VSS.n5121 VSS.n457 258.334
R2396 VSS.n5103 VSS.n488 258.334
R2397 VSS.n4525 VSS.n4524 258.334
R2398 VSS.n4396 VSS.n4395 258.334
R2399 VSS.n4360 VSS.n1750 258.334
R2400 VSS.n3605 VSS.n3487 258.334
R2401 VSS.n4495 VSS.n1474 258.334
R2402 VSS.n4477 VSS.n1508 258.334
R2403 VSS.n4888 VSS.n4887 258.334
R2404 VSS.n4868 VSS.n995 258.334
R2405 VSS.n4850 VSS.n1029 258.334
R2406 VSS.n2078 VSS.n263 258.334
R2407 VSS.n2737 VSS.n2736 258.334
R2408 VSS.n2855 VSS.n512 258.334
R2409 VSS.n3043 VSS.n3042 258.334
R2410 VSS.n3278 VSS.n1532 258.334
R2411 VSS.n3951 VSS.n3950 258.334
R2412 VSS.n2658 VSS.n2657 258.334
R2413 VSS.n2622 VSS.n2621 254.34
R2414 VSS.n2683 VSS.n2582 254.34
R2415 VSS.n2387 VSS.n267 254.34
R2416 VSS.n2267 VSS.n2264 254.34
R2417 VSS.n2299 VSS.n2297 254.34
R2418 VSS.n4159 VSS.n4158 254.34
R2419 VSS.n4212 VSS.n1851 254.34
R2420 VSS.n2542 VSS.n2516 254.34
R2421 VSS.n1883 VSS 252.274
R2422 VSS.n1897 VSS.n1896 251.118
R2423 VSS.n2435 VSS.n1794 250
R2424 VSS.n4146 VSS.n1816 250
R2425 VSS.n3218 VSS.n1930 250
R2426 VSS.n1977 VSS.n1096 250
R2427 VSS.n3056 VSS.n2002 250
R2428 VSS.n3828 VSS.n1039 250
R2429 VSS.n3415 VSS.n3414 250
R2430 VSS.n533 VSS.n532 250
R2431 VSS.n565 VSS.n108 250
R2432 VSS.n630 VSS.n629 250
R2433 VSS.n889 VSS.n407 250
R2434 VSS.n892 VSS.n891 250
R2435 VSS.n5529 VSS.n30 250
R2436 VSS.n3495 VSS.n3491 250
R2437 VSS.n1586 VSS.n1585 250
R2438 VSS.n3447 VSS.n822 250
R2439 VSS.n3803 VSS.n3802 250
R2440 VSS.n2204 VSS.n249 250
R2441 VSS.n2170 VSS.n2168 250
R2442 VSS.n2983 VSS.n498 250
R2443 VSS.n2949 VSS.n2947 250
R2444 VSS.n3380 VSS.n1518 250
R2445 VSS.n3346 VSS.n3344 250
R2446 VSS.n2750 VSS.n2045 250
R2447 VSS.n2624 VSS.n2590 249.663
R2448 VSS.n4627 VSS.n1400 243.201
R2449 VSS.n4660 VSS.n4659 243.201
R2450 VSS.n97 VSS.t42 240.257
R2451 VSS.n396 VSS.t42 240.257
R2452 VSS.n811 VSS.t42 240.257
R2453 VSS.n5474 VSS.t42 240.257
R2454 VSS.n4624 VSS.n4621 236.8
R2455 VSS.n4662 VSS.n4661 236.8
R2456 VSS.n5424 VSS.t42 235.547
R2457 VSS.n5211 VSS.t42 235.547
R2458 VSS.n4958 VSS.t42 235.547
R2459 VSS.n5472 VSS.t42 235.547
R2460 VSS.n1890 VSS.n1889 234
R2461 VSS.t8 VSS.n2544 229.212
R2462 VSS.n1875 VSS.t19 228.745
R2463 VSS.n1877 VSS.t84 228.215
R2464 VSS.n1876 VSS.t86 228.215
R2465 VSS.n1875 VSS.t80 228.215
R2466 VSS.n4282 VSS.n4281 221.667
R2467 VSS.t42 VSS.n128 221.413
R2468 VSS.n5166 VSS.t42 221.413
R2469 VSS.n4913 VSS.t42 221.413
R2470 VSS.n3630 VSS.t42 221.413
R2471 VSS.t42 VSS.n14 221.413
R2472 VSS.t85 VSS.n1883 213.636
R2473 VSS.n1878 VSS.t68 212.96
R2474 VSS.n1893 VSS.t36 212.959
R2475 VSS.n2546 VSS.n2545 212.281
R2476 VSS.t38 VSS.n2627 207.214
R2477 VSS.t38 VSS.n2796 207.214
R2478 VSS.t38 VSS.n3130 207.214
R2479 VSS.t38 VSS.n3188 207.214
R2480 VSS.n4106 VSS.t38 207.214
R2481 VSS.n5398 VSS.t42 202.571
R2482 VSS.n5185 VSS.t42 202.571
R2483 VSS.n4932 VSS.t42 202.571
R2484 VSS.n3654 VSS.t42 202.571
R2485 VSS.t42 VSS.n15 202.571
R2486 VSS.n4629 VSS.n4628 201.927
R2487 VSS.n5562 VSS.n5 197
R2488 VSS.n4677 VSS.n4676 192.796
R2489 VSS.n4676 VSS.n4675 192.796
R2490 VSS.n4675 VSS.n1363 192.796
R2491 VSS.n4669 VSS.n1363 192.796
R2492 VSS.n4669 VSS.n4668 192.796
R2493 VSS.n2525 VSS.n1368 192.796
R2494 VSS.n2526 VSS.n2525 192.796
R2495 VSS.n2528 VSS.n2526 192.796
R2496 VSS.n2528 VSS.n2527 192.796
R2497 VSS.n2527 VSS.n2390 192.796
R2498 VSS.n2544 VSS.n2391 192.796
R2499 VSS.n2539 VSS.n2391 192.796
R2500 VSS.n2539 VSS.n2538 192.796
R2501 VSS.n2538 VSS.n2537 192.796
R2502 VSS.n2537 VSS.n2533 192.796
R2503 VSS.n4656 VSS.n1379 192.796
R2504 VSS.n4650 VSS.n1379 192.796
R2505 VSS.n4650 VSS.n4649 192.796
R2506 VSS.n4649 VSS.n4648 192.796
R2507 VSS.n4648 VSS.n1385 192.796
R2508 VSS.n4642 VSS.n1385 192.796
R2509 VSS.n1403 VSS.n1392 192.796
R2510 VSS.n4616 VSS.n1404 192.796
R2511 VSS.n4610 VSS.n1404 192.796
R2512 VSS.n4608 VSS.n4607 192.796
R2513 VSS.n4607 VSS.n4606 192.796
R2514 VSS.n4606 VSS.n4592 192.796
R2515 VSS.n4600 VSS.n4592 192.796
R2516 VSS.n4600 VSS.n4599 192.796
R2517 VSS.n4599 VSS.n4598 192.796
R2518 VSS.n5540 VSS.n5539 192.796
R2519 VSS.n5541 VSS.n5540 192.796
R2520 VSS.n5541 VSS.n16 192.796
R2521 VSS.n5547 VSS.n16 192.796
R2522 VSS.n5548 VSS.n5547 192.796
R2523 VSS.n5549 VSS.n9 192.796
R2524 VSS.n5556 VSS.n9 192.796
R2525 VSS.n5557 VSS.n5556 192.796
R2526 VSS.n5558 VSS.n5557 192.796
R2527 VSS.n5558 VSS.n4 192.796
R2528 VSS.n5563 VSS.n4 192.796
R2529 VSS.n2642 VSS.t38 189.579
R2530 VSS.n2811 VSS.t38 189.579
R2531 VSS.n3132 VSS.t38 189.579
R2532 VSS.n3234 VSS.t38 189.579
R2533 VSS.n4120 VSS.t38 189.579
R2534 VSS.n5372 VSS.n5369 187.249
R2535 VSS.n2609 VSS.t38 186.55
R2536 VSS.t33 VSS.n1180 186.55
R2537 VSS.n2557 VSS.t31 186.55
R2538 VSS.n2376 VSS.t40 186.55
R2539 VSS.n2312 VSS.t44 186.55
R2540 VSS.t42 VSS.n5385 186.55
R2541 VSS.n2452 VSS.n2451 185
R2542 VSS.n2450 VSS.n2449 185
R2543 VSS.n2448 VSS.n2447 185
R2544 VSS.n2446 VSS.n2445 185
R2545 VSS.n2444 VSS.n2443 185
R2546 VSS.n2442 VSS.n2441 185
R2547 VSS.n2440 VSS.n2439 185
R2548 VSS.n2438 VSS.n2437 185
R2549 VSS.n2436 VSS.n2435 185
R2550 VSS.n4131 VSS.n4130 185
R2551 VSS.n4133 VSS.n4132 185
R2552 VSS.n4135 VSS.n4134 185
R2553 VSS.n4137 VSS.n4136 185
R2554 VSS.n4139 VSS.n4138 185
R2555 VSS.n4141 VSS.n4140 185
R2556 VSS.n4143 VSS.n4142 185
R2557 VSS.n4145 VSS.n4144 185
R2558 VSS.n4147 VSS.n4146 185
R2559 VSS.n4095 VSS.n4094 185
R2560 VSS.n4093 VSS.n4092 185
R2561 VSS.n4091 VSS.n4090 185
R2562 VSS.n4089 VSS.n4088 185
R2563 VSS.n4087 VSS.n4086 185
R2564 VSS.n4085 VSS.n4084 185
R2565 VSS.n4083 VSS.n4082 185
R2566 VSS.n1832 VSS.n1831 185
R2567 VSS.n4275 VSS.n4274 185
R2568 VSS.n3203 VSS.n1926 185
R2569 VSS.n3205 VSS.n3204 185
R2570 VSS.n3207 VSS.n3206 185
R2571 VSS.n3209 VSS.n3208 185
R2572 VSS.n3211 VSS.n3210 185
R2573 VSS.n3213 VSS.n3212 185
R2574 VSS.n3215 VSS.n3214 185
R2575 VSS.n3217 VSS.n3216 185
R2576 VSS.n3219 VSS.n3218 185
R2577 VSS.n3251 VSS.n3250 185
R2578 VSS.n3253 VSS.n3252 185
R2579 VSS.n3255 VSS.n3254 185
R2580 VSS.n3257 VSS.n3256 185
R2581 VSS.n3259 VSS.n3258 185
R2582 VSS.n3261 VSS.n3260 185
R2583 VSS.n3263 VSS.n3262 185
R2584 VSS.n3265 VSS.n3264 185
R2585 VSS.n3266 VSS.n1944 185
R2586 VSS.n1962 VSS.n1961 185
R2587 VSS.n1964 VSS.n1963 185
R2588 VSS.n1966 VSS.n1965 185
R2589 VSS.n1968 VSS.n1967 185
R2590 VSS.n1970 VSS.n1969 185
R2591 VSS.n1972 VSS.n1971 185
R2592 VSS.n1974 VSS.n1973 185
R2593 VSS.n1976 VSS.n1975 185
R2594 VSS.n1978 VSS.n1977 185
R2595 VSS.n3109 VSS.n3108 185
R2596 VSS.n3106 VSS.n3105 185
R2597 VSS.n3104 VSS.n3103 185
R2598 VSS.n3102 VSS.n3101 185
R2599 VSS.n3100 VSS.n3099 185
R2600 VSS.n1112 VSS.n1111 185
R2601 VSS.n4773 VSS.n4772 185
R2602 VSS.n4771 VSS.n1110 185
R2603 VSS.n4770 VSS.n4769 185
R2604 VSS.n2899 VSS.n2898 185
R2605 VSS.n2897 VSS.n2896 185
R2606 VSS.n2895 VSS.n2894 185
R2607 VSS.n2893 VSS.n2892 185
R2608 VSS.n2891 VSS.n2890 185
R2609 VSS.n2889 VSS.n2888 185
R2610 VSS.n2887 VSS.n2886 185
R2611 VSS.n2885 VSS.n2884 185
R2612 VSS.n2883 VSS.n2002 185
R2613 VSS.n2828 VSS.n2827 185
R2614 VSS.n2830 VSS.n2829 185
R2615 VSS.n2832 VSS.n2831 185
R2616 VSS.n2834 VSS.n2833 185
R2617 VSS.n2836 VSS.n2835 185
R2618 VSS.n2838 VSS.n2837 185
R2619 VSS.n2840 VSS.n2839 185
R2620 VSS.n2842 VSS.n2841 185
R2621 VSS.n2843 VSS.n2020 185
R2622 VSS.n4793 VSS.n1053 185
R2623 VSS.n4844 VSS.n4843 185
R2624 VSS.n4842 VSS.n1054 185
R2625 VSS.n4841 VSS.n4840 185
R2626 VSS.n4839 VSS.n4838 185
R2627 VSS.n4837 VSS.n4836 185
R2628 VSS.n4835 VSS.n4834 185
R2629 VSS.n4833 VSS.n4832 185
R2630 VSS.n4831 VSS.n4830 185
R2631 VSS.n1128 VSS.n1086 185
R2632 VSS.n1127 VSS.n1126 185
R2633 VSS.n1125 VSS.n1124 185
R2634 VSS.n1123 VSS.n1122 185
R2635 VSS.n1121 VSS.n1120 185
R2636 VSS.n1119 VSS.n1118 185
R2637 VSS.n1117 VSS.n1116 185
R2638 VSS.n1115 VSS.n1114 185
R2639 VSS.n1113 VSS.n1055 185
R2640 VSS.n3432 VSS.n3431 185
R2641 VSS.n3430 VSS.n3429 185
R2642 VSS.n3428 VSS.n3427 185
R2643 VSS.n3426 VSS.n3425 185
R2644 VSS.n3424 VSS.n3423 185
R2645 VSS.n3422 VSS.n3421 185
R2646 VSS.n3420 VSS.n3419 185
R2647 VSS.n3418 VSS.n3417 185
R2648 VSS.n3416 VSS.n3415 185
R2649 VSS.n3813 VSS.n3812 185
R2650 VSS.n3815 VSS.n3814 185
R2651 VSS.n3817 VSS.n3816 185
R2652 VSS.n3819 VSS.n3818 185
R2653 VSS.n3821 VSS.n3820 185
R2654 VSS.n3823 VSS.n3822 185
R2655 VSS.n3825 VSS.n3824 185
R2656 VSS.n3827 VSS.n3826 185
R2657 VSS.n3829 VSS.n3828 185
R2658 VSS.n266 VSS.n239 185
R2659 VSS.n2341 VSS.n2340 185
R2660 VSS.n2343 VSS.n2342 185
R2661 VSS.n2345 VSS.n2344 185
R2662 VSS.n2347 VSS.n2346 185
R2663 VSS.n2349 VSS.n2348 185
R2664 VSS.n2351 VSS.n2350 185
R2665 VSS.n2353 VSS.n2352 185
R2666 VSS.n2355 VSS.n2354 185
R2667 VSS.n550 VSS.n549 185
R2668 VSS.n548 VSS.n547 185
R2669 VSS.n546 VSS.n545 185
R2670 VSS.n544 VSS.n543 185
R2671 VSS.n542 VSS.n541 185
R2672 VSS.n540 VSS.n539 185
R2673 VSS.n538 VSS.n537 185
R2674 VSS.n536 VSS.n535 185
R2675 VSS.n534 VSS.n533 185
R2676 VSS.n5352 VSS.n5351 185
R2677 VSS.n5354 VSS.n5353 185
R2678 VSS.n5356 VSS.n5355 185
R2679 VSS.n5358 VSS.n5357 185
R2680 VSS.n5360 VSS.n5359 185
R2681 VSS.n5362 VSS.n5361 185
R2682 VSS.n5364 VSS.n5363 185
R2683 VSS.n5366 VSS.n5365 185
R2684 VSS.n5367 VSS.n122 185
R2685 VSS.n2339 VSS.n200 185
R2686 VSS.n2338 VSS.n2337 185
R2687 VSS.n2336 VSS.n2335 185
R2688 VSS.n2334 VSS.n2333 185
R2689 VSS.n2332 VSS.n2331 185
R2690 VSS.n2330 VSS.n2329 185
R2691 VSS.n2328 VSS.n2327 185
R2692 VSS.n2326 VSS.n2325 185
R2693 VSS.n2324 VSS.n2323 185
R2694 VSS.n597 VSS.n596 185
R2695 VSS.n599 VSS.n598 185
R2696 VSS.n601 VSS.n600 185
R2697 VSS.n603 VSS.n602 185
R2698 VSS.n605 VSS.n604 185
R2699 VSS.n607 VSS.n606 185
R2700 VSS.n609 VSS.n608 185
R2701 VSS.n611 VSS.n610 185
R2702 VSS.n629 VSS.n612 185
R2703 VSS.n104 VSS.n101 185
R2704 VSS.n552 VSS.n551 185
R2705 VSS.n554 VSS.n553 185
R2706 VSS.n556 VSS.n555 185
R2707 VSS.n558 VSS.n557 185
R2708 VSS.n560 VSS.n559 185
R2709 VSS.n562 VSS.n561 185
R2710 VSS.n564 VSS.n563 185
R2711 VSS.n566 VSS.n565 185
R2712 VSS.n588 VSS.n108 185
R2713 VSS.t41 VSS.n108 185
R2714 VSS.n586 VSS.n585 185
R2715 VSS.n579 VSS.n578 185
R2716 VSS.n577 VSS.n576 185
R2717 VSS.n5337 VSS.n5336 185
R2718 VSS.n5335 VSS.n5334 185
R2719 VSS.n176 VSS.n175 185
R2720 VSS.n174 VSS.n173 185
R2721 VSS.n5350 VSS.n5349 185
R2722 VSS.n568 VSS.n567 185
R2723 VSS.n587 VSS.n190 185
R2724 VSS.t72 VSS.n190 185
R2725 VSS.n571 VSS.n570 185
R2726 VSS.n573 VSS.n181 185
R2727 VSS.n5333 VSS.n5332 185
R2728 VSS.n184 VSS.n180 185
R2729 VSS.n183 VSS.n182 185
R2730 VSS.n5346 VSS.n5345 185
R2731 VSS.n5348 VSS.n5347 185
R2732 VSS.n631 VSS.n630 185
R2733 VSS.n627 VSS.n626 185
R2734 VSS.n625 VSS.n624 185
R2735 VSS.n5315 VSS.n5314 185
R2736 VSS.n5317 VSS.n5316 185
R2737 VSS.n215 VSS.n214 185
R2738 VSS.n213 VSS.n207 185
R2739 VSS.n206 VSS.n201 185
R2740 VSS.n5330 VSS.n5329 185
R2741 VSS.t72 VSS.n5330 185
R2742 VSS.n614 VSS.n613 185
R2743 VSS.n628 VSS.n229 185
R2744 VSS.t39 VSS.n229 185
R2745 VSS.n623 VSS.n220 185
R2746 VSS.n5313 VSS.n5312 185
R2747 VSS.n219 VSS.n217 185
R2748 VSS.n225 VSS.n216 185
R2749 VSS.n224 VSS.n223 185
R2750 VSS.n5326 VSS.n5325 185
R2751 VSS.n5328 VSS.n5327 185
R2752 VSS.n403 VSS.n400 185
R2753 VSS.n876 VSS.n875 185
R2754 VSS.n878 VSS.n877 185
R2755 VSS.n880 VSS.n879 185
R2756 VSS.n882 VSS.n881 185
R2757 VSS.n884 VSS.n883 185
R2758 VSS.n886 VSS.n885 185
R2759 VSS.n888 VSS.n887 185
R2760 VSS.n890 VSS.n889 185
R2761 VSS.n531 VSS.n457 185
R2762 VSS.n530 VSS.n529 185
R2763 VSS.n528 VSS.n527 185
R2764 VSS.n526 VSS.n525 185
R2765 VSS.n524 VSS.n523 185
R2766 VSS.n522 VSS.n521 185
R2767 VSS.n520 VSS.n519 185
R2768 VSS.n518 VSS.n517 185
R2769 VSS.n516 VSS.n515 185
R2770 VSS.n5142 VSS.n5141 185
R2771 VSS.n5144 VSS.n5143 185
R2772 VSS.n5146 VSS.n5145 185
R2773 VSS.n5148 VSS.n5147 185
R2774 VSS.n5150 VSS.n5149 185
R2775 VSS.n5152 VSS.n5151 185
R2776 VSS.n5154 VSS.n5153 185
R2777 VSS.n5156 VSS.n5155 185
R2778 VSS.n5157 VSS.n421 185
R2779 VSS.n873 VSS.n407 185
R2780 VSS.t53 VSS.n407 185
R2781 VSS.n867 VSS.n866 185
R2782 VSS.n862 VSS.n861 185
R2783 VSS.n860 VSS.n859 185
R2784 VSS.n5127 VSS.n5126 185
R2785 VSS.n5129 VSS.n5128 185
R2786 VSS.n430 VSS.n429 185
R2787 VSS.n428 VSS.n427 185
R2788 VSS.n5140 VSS.n5139 185
R2789 VSS.n958 VSS.n874 185
R2790 VSS.n863 VSS.n849 185
R2791 VSS.n865 VSS.n864 185
R2792 VSS.n858 VSS.n439 185
R2793 VSS.n5125 VSS.n5124 185
R2794 VSS.n441 VSS.n437 185
R2795 VSS.n440 VSS.n436 185
R2796 VSS.n5136 VSS.n5135 185
R2797 VSS.n5138 VSS.n5137 185
R2798 VSS.n697 VSS.n488 185
R2799 VSS.n696 VSS.n695 185
R2800 VSS.n694 VSS.n693 185
R2801 VSS.n692 VSS.n691 185
R2802 VSS.n690 VSS.n689 185
R2803 VSS.n688 VSS.n687 185
R2804 VSS.n686 VSS.n685 185
R2805 VSS.n684 VSS.n683 185
R2806 VSS.n682 VSS.n681 185
R2807 VSS.n909 VSS.n908 185
R2808 VSS.n907 VSS.n906 185
R2809 VSS.n905 VSS.n904 185
R2810 VSS.n903 VSS.n902 185
R2811 VSS.n901 VSS.n900 185
R2812 VSS.n899 VSS.n898 185
R2813 VSS.n897 VSS.n896 185
R2814 VSS.n895 VSS.n894 185
R2815 VSS.n893 VSS.n892 185
R2816 VSS.n960 VSS.n959 185
R2817 VSS.n957 VSS.n956 185
R2818 VSS.n955 VSS.n954 185
R2819 VSS.n953 VSS.n952 185
R2820 VSS.n951 VSS.n950 185
R2821 VSS.n949 VSS.n948 185
R2822 VSS.n947 VSS.n946 185
R2823 VSS.n945 VSS.n944 185
R2824 VSS.n943 VSS.n942 185
R2825 VSS.n4524 VSS.n4507 185
R2826 VSS.n4522 VSS.n4521 185
R2827 VSS.n4520 VSS.n4508 185
R2828 VSS.n4519 VSS.n4518 185
R2829 VSS.n4516 VSS.n4509 185
R2830 VSS.n4514 VSS.n4513 185
R2831 VSS.n4512 VSS.n4511 185
R2832 VSS.n56 VSS.n55 185
R2833 VSS.n5481 VSS.n5480 185
R2834 VSS.n4314 VSS.n1750 185
R2835 VSS.n4313 VSS.n4312 185
R2836 VSS.n4311 VSS.n4310 185
R2837 VSS.n4309 VSS.n4308 185
R2838 VSS.n4307 VSS.n4306 185
R2839 VSS.n4305 VSS.n4304 185
R2840 VSS.n4303 VSS.n4302 185
R2841 VSS.n4301 VSS.n4300 185
R2842 VSS.n4299 VSS.n4298 185
R2843 VSS.n4395 VSS.n4394 185
R2844 VSS.n4393 VSS.n4392 185
R2845 VSS.n4391 VSS.n4390 185
R2846 VSS.n4389 VSS.n4388 185
R2847 VSS.n4387 VSS.n4386 185
R2848 VSS.n4385 VSS.n4384 185
R2849 VSS.n4383 VSS.n4382 185
R2850 VSS.n4381 VSS.n4380 185
R2851 VSS.n1450 VSS.n1442 185
R2852 VSS.n1736 VSS.n1411 185
R2853 VSS.n1727 VSS.n1726 185
R2854 VSS.n1722 VSS.n1721 185
R2855 VSS.n1720 VSS.n1719 185
R2856 VSS.n4368 VSS.n4367 185
R2857 VSS.n4366 VSS.n4365 185
R2858 VSS.n1696 VSS.n1695 185
R2859 VSS.n1694 VSS.n1693 185
R2860 VSS.n4397 VSS.n4396 185
R2861 VSS.n1738 VSS.n1737 185
R2862 VSS.n1723 VSS.n1711 185
R2863 VSS.n1725 VSS.n1724 185
R2864 VSS.n1718 VSS.n1702 185
R2865 VSS.n4364 VSS.n4363 185
R2866 VSS.n1705 VSS.n1701 185
R2867 VSS.n1704 VSS.n1703 185
R2868 VSS.n4377 VSS.n4376 185
R2869 VSS.n4379 VSS.n4378 185
R2870 VSS.n1434 VSS.n28 185
R2871 VSS.n1432 VSS.n1431 185
R2872 VSS.n1430 VSS.n1421 185
R2873 VSS.n1429 VSS.n1428 185
R2874 VSS.n1427 VSS.n1426 185
R2875 VSS.n1425 VSS.n1424 185
R2876 VSS.n1423 VSS.n1422 185
R2877 VSS.n1410 VSS.n1409 185
R2878 VSS.n4582 VSS.n4581 185
R2879 VSS.n5515 VSS.n35 185
R2880 VSS.n5517 VSS.n5516 185
R2881 VSS.n5519 VSS.n33 185
R2882 VSS.n5521 VSS.n5520 185
R2883 VSS.n5522 VSS.n32 185
R2884 VSS.n5524 VSS.n5523 185
R2885 VSS.n5526 VSS.n31 185
R2886 VSS.n5527 VSS.n29 185
R2887 VSS.n5530 VSS.n5529 185
R2888 VSS.n4544 VSS.n30 185
R2889 VSS.t56 VSS.n30 185
R2890 VSS.n4553 VSS.n4552 185
R2891 VSS.n4556 VSS.n4555 185
R2892 VSS.n4542 VSS.n4540 185
R2893 VSS.n4530 VSS.n4528 185
R2894 VSS.n4568 VSS.n4567 185
R2895 VSS.n4571 VSS.n4570 185
R2896 VSS.n4527 VSS.n1445 185
R2897 VSS.n4525 VSS.n1444 185
R2898 VSS.n1433 VSS.n27 185
R2899 VSS.n4551 VSS.n4550 185
R2900 VSS.n4549 VSS.n4539 185
R2901 VSS.n4538 VSS.n4537 185
R2902 VSS.n4536 VSS.n4535 185
R2903 VSS.n4566 VSS.n4565 185
R2904 VSS.n4564 VSS.n1449 185
R2905 VSS.n1448 VSS.n1443 185
R2906 VSS.n4578 VSS.n4577 185
R2907 VSS.n3512 VSS.n3511 185
R2908 VSS.n3510 VSS.n3497 185
R2909 VSS.n3509 VSS.n3508 185
R2910 VSS.n3507 VSS.n3506 185
R2911 VSS.n3505 VSS.n3504 185
R2912 VSS.n3503 VSS.n3502 185
R2913 VSS.n3501 VSS.n3500 185
R2914 VSS.n3499 VSS.n3498 185
R2915 VSS.n3495 VSS.n1452 185
R2916 VSS.n3587 VSS.n1474 185
R2917 VSS.n3589 VSS.n3588 185
R2918 VSS.n3591 VSS.n3590 185
R2919 VSS.n3593 VSS.n3592 185
R2920 VSS.n3595 VSS.n3594 185
R2921 VSS.n3597 VSS.n3596 185
R2922 VSS.n3599 VSS.n3598 185
R2923 VSS.n3601 VSS.n3600 185
R2924 VSS.n3603 VSS.n3602 185
R2925 VSS.n3606 VSS.n3605 185
R2926 VSS.n3608 VSS.n3607 185
R2927 VSS.n3610 VSS.n3609 185
R2928 VSS.n3612 VSS.n3611 185
R2929 VSS.n3614 VSS.n3613 185
R2930 VSS.n3616 VSS.n3615 185
R2931 VSS.n3618 VSS.n3617 185
R2932 VSS.n3620 VSS.n3619 185
R2933 VSS.n3621 VSS.n3569 185
R2934 VSS.n3539 VSS.n3491 185
R2935 VSS.t54 VSS.n3491 185
R2936 VSS.n3548 VSS.n3547 185
R2937 VSS.n3536 VSS.n3516 185
R2938 VSS.n3561 VSS.n3560 185
R2939 VSS.n3518 VSS.n3515 185
R2940 VSS.n3521 VSS.n3520 185
R2941 VSS.n3522 VSS.n3485 185
R2942 VSS.n3673 VSS.n3672 185
R2943 VSS.n3487 VSS.n3486 185
R2944 VSS.n4498 VSS.n1456 185
R2945 VSS.n3546 VSS.n1457 185
R2946 VSS.n3538 VSS.n3537 185
R2947 VSS.n3559 VSS.n3558 185
R2948 VSS.n3557 VSS.n3556 185
R2949 VSS.n3531 VSS.n3530 185
R2950 VSS.n3529 VSS.n3528 185
R2951 VSS.n3484 VSS.n3483 185
R2952 VSS.n3482 VSS.n3481 185
R2953 VSS.n1535 VSS.n1508 185
R2954 VSS.n3571 VSS.n3570 185
R2955 VSS.n3573 VSS.n3572 185
R2956 VSS.n3575 VSS.n3574 185
R2957 VSS.n3577 VSS.n3576 185
R2958 VSS.n3579 VSS.n3578 185
R2959 VSS.n3581 VSS.n3580 185
R2960 VSS.n3583 VSS.n3582 185
R2961 VSS.n3585 VSS.n3584 185
R2962 VSS.n1603 VSS.n1602 185
R2963 VSS.n1601 VSS.n1600 185
R2964 VSS.n1599 VSS.n1598 185
R2965 VSS.n1597 VSS.n1596 185
R2966 VSS.n1595 VSS.n1594 185
R2967 VSS.n1593 VSS.n1592 185
R2968 VSS.n1591 VSS.n1590 185
R2969 VSS.n1589 VSS.n1588 185
R2970 VSS.n1587 VSS.n1586 185
R2971 VSS.n4500 VSS.n4499 185
R2972 VSS.n1604 VSS.n1454 185
R2973 VSS.n1606 VSS.n1605 185
R2974 VSS.n1608 VSS.n1607 185
R2975 VSS.n1610 VSS.n1609 185
R2976 VSS.n1612 VSS.n1611 185
R2977 VSS.n1614 VSS.n1613 185
R2978 VSS.n1616 VSS.n1615 185
R2979 VSS.n1618 VSS.n1617 185
R2980 VSS.n1643 VSS.n1642 185
R2981 VSS.n1641 VSS.n1640 185
R2982 VSS.n1634 VSS.n1633 185
R2983 VSS.n1632 VSS.n1631 185
R2984 VSS.n4482 VSS.n4481 185
R2985 VSS.n4484 VSS.n4483 185
R2986 VSS.n1481 VSS.n1480 185
R2987 VSS.n1479 VSS.n1473 185
R2988 VSS.n4495 VSS.n4494 185
R2989 VSS.n1620 VSS.n1619 185
R2990 VSS.n1622 VSS.n1498 185
R2991 VSS.t49 VSS.n1498 185
R2992 VSS.n1624 VSS.n1623 185
R2993 VSS.n1626 VSS.n1490 185
R2994 VSS.n4480 VSS.n4479 185
R2995 VSS.n1492 VSS.n1488 185
R2996 VSS.n1491 VSS.n1487 185
R2997 VSS.n4491 VSS.n4490 185
R2998 VSS.n4493 VSS.n4492 185
R2999 VSS.n818 VSS.n815 185
R3000 VSS.n3434 VSS.n3433 185
R3001 VSS.n3436 VSS.n3435 185
R3002 VSS.n3438 VSS.n3437 185
R3003 VSS.n3440 VSS.n3439 185
R3004 VSS.n3442 VSS.n3441 185
R3005 VSS.n3444 VSS.n3443 185
R3006 VSS.n3446 VSS.n3445 185
R3007 VSS.n3448 VSS.n3447 185
R3008 VSS.n4810 VSS.n995 185
R3009 VSS.n4809 VSS.n4808 185
R3010 VSS.n4807 VSS.n4806 185
R3011 VSS.n4805 VSS.n4804 185
R3012 VSS.n4803 VSS.n4802 185
R3013 VSS.n4801 VSS.n4800 185
R3014 VSS.n4799 VSS.n4798 185
R3015 VSS.n4797 VSS.n4796 185
R3016 VSS.n4795 VSS.n4794 185
R3017 VSS.n4889 VSS.n4888 185
R3018 VSS.n4891 VSS.n4890 185
R3019 VSS.n4893 VSS.n4892 185
R3020 VSS.n4895 VSS.n4894 185
R3021 VSS.n4897 VSS.n4896 185
R3022 VSS.n4899 VSS.n4898 185
R3023 VSS.n4901 VSS.n4900 185
R3024 VSS.n4903 VSS.n4902 185
R3025 VSS.n4904 VSS.n836 185
R3026 VSS.n3450 VSS.n822 185
R3027 VSS.t65 VSS.n822 185
R3028 VSS.n3453 VSS.n3452 185
R3029 VSS.n3460 VSS.n3454 185
R3030 VSS.n3462 VSS.n3461 185
R3031 VSS.n4874 VSS.n4873 185
R3032 VSS.n4876 VSS.n4875 185
R3033 VSS.n845 VSS.n844 185
R3034 VSS.n843 VSS.n842 185
R3035 VSS.n4887 VSS.n4886 185
R3036 VSS.n3686 VSS.n3685 185
R3037 VSS.n3472 VSS.n3471 185
R3038 VSS.n3470 VSS.n3469 185
R3039 VSS.n3463 VSS.n977 185
R3040 VSS.n4872 VSS.n4871 185
R3041 VSS.n979 VSS.n975 185
R3042 VSS.n978 VSS.n974 185
R3043 VSS.n4883 VSS.n4882 185
R3044 VSS.n4885 VSS.n4884 185
R3045 VSS.n4828 VSS.n1029 185
R3046 VSS.n4827 VSS.n4826 185
R3047 VSS.n4825 VSS.n4824 185
R3048 VSS.n4823 VSS.n4822 185
R3049 VSS.n4821 VSS.n4820 185
R3050 VSS.n4819 VSS.n4818 185
R3051 VSS.n4817 VSS.n4816 185
R3052 VSS.n4815 VSS.n4814 185
R3053 VSS.n4813 VSS.n4812 185
R3054 VSS.n3738 VSS.n3737 185
R3055 VSS.n3740 VSS.n3739 185
R3056 VSS.n3742 VSS.n3741 185
R3057 VSS.n3744 VSS.n3743 185
R3058 VSS.n3746 VSS.n3745 185
R3059 VSS.n3748 VSS.n3747 185
R3060 VSS.n3750 VSS.n3749 185
R3061 VSS.n3752 VSS.n3751 185
R3062 VSS.n3802 VSS.n3753 185
R3063 VSS.n3688 VSS.n3687 185
R3064 VSS.n3690 VSS.n3689 185
R3065 VSS.n3692 VSS.n3691 185
R3066 VSS.n3694 VSS.n3693 185
R3067 VSS.n3696 VSS.n3695 185
R3068 VSS.n3698 VSS.n3697 185
R3069 VSS.n3700 VSS.n3699 185
R3070 VSS.n3702 VSS.n3701 185
R3071 VSS.n3704 VSS.n3703 185
R3072 VSS.n3729 VSS.n3728 185
R3073 VSS.n3727 VSS.n3726 185
R3074 VSS.n3720 VSS.n3719 185
R3075 VSS.n3718 VSS.n3717 185
R3076 VSS.n4855 VSS.n4854 185
R3077 VSS.n4857 VSS.n4856 185
R3078 VSS.n1002 VSS.n1001 185
R3079 VSS.n1000 VSS.n994 185
R3080 VSS.n4868 VSS.n4867 185
R3081 VSS.n3706 VSS.n3705 185
R3082 VSS.n3708 VSS.n1019 185
R3083 VSS.t69 VSS.n1019 185
R3084 VSS.n3710 VSS.n3709 185
R3085 VSS.n3712 VSS.n1011 185
R3086 VSS.n4853 VSS.n4852 185
R3087 VSS.n1013 VSS.n1009 185
R3088 VSS.n1012 VSS.n1008 185
R3089 VSS.n4864 VSS.n4863 185
R3090 VSS.n4866 VSS.n4865 185
R3091 VSS.n934 VSS.n933 185
R3092 VSS.n932 VSS.n931 185
R3093 VSS.n925 VSS.n924 185
R3094 VSS.n923 VSS.n922 185
R3095 VSS.n5108 VSS.n5107 185
R3096 VSS.n5110 VSS.n5109 185
R3097 VSS.n464 VSS.n463 185
R3098 VSS.n462 VSS.n456 185
R3099 VSS.n5121 VSS.n5120 185
R3100 VSS.n911 VSS.n910 185
R3101 VSS.n913 VSS.n478 185
R3102 VSS.t73 VSS.n478 185
R3103 VSS.n915 VSS.n914 185
R3104 VSS.n917 VSS.n470 185
R3105 VSS.n5106 VSS.n5105 185
R3106 VSS.n472 VSS.n468 185
R3107 VSS.n471 VSS.n467 185
R3108 VSS.n5117 VSS.n5116 185
R3109 VSS.n5119 VSS.n5118 185
R3110 VSS.n265 VSS.n263 185
R3111 VSS.n5304 VSS.n5303 185
R3112 VSS.n5302 VSS.n264 185
R3113 VSS.n5301 VSS.n5300 185
R3114 VSS.n5299 VSS.n5298 185
R3115 VSS.n5297 VSS.n5296 185
R3116 VSS.n5295 VSS.n5294 185
R3117 VSS.n5293 VSS.n5292 185
R3118 VSS.n5291 VSS.n5290 185
R3119 VSS.n2736 VSS.n2072 185
R3120 VSS.n2734 VSS.n2733 185
R3121 VSS.n2732 VSS.n2073 185
R3122 VSS.n2731 VSS.n2730 185
R3123 VSS.n2728 VSS.n2074 185
R3124 VSS.n2726 VSS.n2725 185
R3125 VSS.n2724 VSS.n2075 185
R3126 VSS.n2723 VSS.n2722 185
R3127 VSS.n2720 VSS.n2076 185
R3128 VSS.n2187 VSS.n2186 185
R3129 VSS.n2184 VSS.n2100 185
R3130 VSS.n2182 VSS.n2181 185
R3131 VSS.n2180 VSS.n2101 185
R3132 VSS.n2179 VSS.n2178 185
R3133 VSS.n2176 VSS.n2102 185
R3134 VSS.n2174 VSS.n2173 185
R3135 VSS.n2172 VSS.n2103 185
R3136 VSS.n2171 VSS.n2170 185
R3137 VSS.n2189 VSS.n2188 185
R3138 VSS.n2191 VSS.n2190 185
R3139 VSS.n2193 VSS.n2192 185
R3140 VSS.n2195 VSS.n2194 185
R3141 VSS.n2197 VSS.n2196 185
R3142 VSS.n2199 VSS.n2198 185
R3143 VSS.n2201 VSS.n2200 185
R3144 VSS.n2203 VSS.n2202 185
R3145 VSS.n2205 VSS.n2204 185
R3146 VSS.n514 VSS.n512 185
R3147 VSS.n5097 VSS.n5096 185
R3148 VSS.n5095 VSS.n513 185
R3149 VSS.n5094 VSS.n5093 185
R3150 VSS.n5092 VSS.n5091 185
R3151 VSS.n5090 VSS.n5089 185
R3152 VSS.n5088 VSS.n5087 185
R3153 VSS.n5086 VSS.n5085 185
R3154 VSS.n5084 VSS.n5083 185
R3155 VSS.n3042 VSS.n2849 185
R3156 VSS.n3040 VSS.n3039 185
R3157 VSS.n3038 VSS.n2850 185
R3158 VSS.n3037 VSS.n3036 185
R3159 VSS.n3034 VSS.n2851 185
R3160 VSS.n3032 VSS.n3031 185
R3161 VSS.n3030 VSS.n2852 185
R3162 VSS.n3029 VSS.n3028 185
R3163 VSS.n3026 VSS.n2853 185
R3164 VSS.n2966 VSS.n2965 185
R3165 VSS.n2963 VSS.n2879 185
R3166 VSS.n2961 VSS.n2960 185
R3167 VSS.n2959 VSS.n2880 185
R3168 VSS.n2958 VSS.n2957 185
R3169 VSS.n2955 VSS.n2881 185
R3170 VSS.n2953 VSS.n2952 185
R3171 VSS.n2951 VSS.n2882 185
R3172 VSS.n2950 VSS.n2949 185
R3173 VSS.n2968 VSS.n2967 185
R3174 VSS.n2970 VSS.n2969 185
R3175 VSS.n2972 VSS.n2971 185
R3176 VSS.n2974 VSS.n2973 185
R3177 VSS.n2976 VSS.n2975 185
R3178 VSS.n2978 VSS.n2977 185
R3179 VSS.n2980 VSS.n2979 185
R3180 VSS.n2982 VSS.n2981 185
R3181 VSS.n2984 VSS.n2983 185
R3182 VSS.n2877 VSS.n498 185
R3183 VSS.t59 VSS.n498 185
R3184 VSS.n2876 VSS.n2875 185
R3185 VSS.n3000 VSS.n2999 185
R3186 VSS.n3002 VSS.n3001 185
R3187 VSS.n2867 VSS.n2866 185
R3188 VSS.n2865 VSS.n2864 185
R3189 VSS.n3014 VSS.n3013 185
R3190 VSS.n3016 VSS.n3015 185
R3191 VSS.n2856 VSS.n2855 185
R3192 VSS.n2878 VSS.n2874 185
R3193 VSS.n2992 VSS.n2991 185
R3194 VSS.n2992 VSS.t52 185
R3195 VSS.n2998 VSS.n2997 185
R3196 VSS.n2995 VSS.n2868 185
R3197 VSS.n2994 VSS.n2993 185
R3198 VSS.n3009 VSS.n3008 185
R3199 VSS.n3012 VSS.n3011 185
R3200 VSS.n2857 VSS.n2854 185
R3201 VSS.n3024 VSS.n3023 185
R3202 VSS.n2209 VSS.n249 185
R3203 VSS.t30 VSS.n249 185
R3204 VSS.n2099 VSS.n2098 185
R3205 VSS.n2222 VSS.n2221 185
R3206 VSS.n2224 VSS.n2223 185
R3207 VSS.n2090 VSS.n2089 185
R3208 VSS.n2088 VSS.n2087 185
R3209 VSS.n2236 VSS.n2235 185
R3210 VSS.n2238 VSS.n2237 185
R3211 VSS.n2079 VSS.n2078 185
R3212 VSS.n2208 VSS.n2097 185
R3213 VSS.n2214 VSS.n2213 185
R3214 VSS.n2214 VSS.t57 185
R3215 VSS.n2220 VSS.n2219 185
R3216 VSS.n2217 VSS.n2091 185
R3217 VSS.n2216 VSS.n2215 185
R3218 VSS.n2231 VSS.n2230 185
R3219 VSS.n2234 VSS.n2233 185
R3220 VSS.n2080 VSS.n2077 185
R3221 VSS.n2718 VSS.n2717 185
R3222 VSS.n1534 VSS.n1532 185
R3223 VSS.n4471 VSS.n4470 185
R3224 VSS.n4469 VSS.n1533 185
R3225 VSS.n4468 VSS.n4467 185
R3226 VSS.n4466 VSS.n4465 185
R3227 VSS.n4464 VSS.n4463 185
R3228 VSS.n4462 VSS.n4461 185
R3229 VSS.n4460 VSS.n4459 185
R3230 VSS.n4458 VSS.n4457 185
R3231 VSS.n3950 VSS.n3272 185
R3232 VSS.n3948 VSS.n3947 185
R3233 VSS.n3946 VSS.n3273 185
R3234 VSS.n3945 VSS.n3944 185
R3235 VSS.n3942 VSS.n3274 185
R3236 VSS.n3940 VSS.n3939 185
R3237 VSS.n3938 VSS.n3275 185
R3238 VSS.n3937 VSS.n3936 185
R3239 VSS.n3934 VSS.n3276 185
R3240 VSS.n3363 VSS.n3362 185
R3241 VSS.n3360 VSS.n3302 185
R3242 VSS.n3358 VSS.n3357 185
R3243 VSS.n3356 VSS.n3303 185
R3244 VSS.n3355 VSS.n3354 185
R3245 VSS.n3352 VSS.n3304 185
R3246 VSS.n3350 VSS.n3349 185
R3247 VSS.n3348 VSS.n3305 185
R3248 VSS.n3347 VSS.n3346 185
R3249 VSS.n3365 VSS.n3364 185
R3250 VSS.n3367 VSS.n3366 185
R3251 VSS.n3369 VSS.n3368 185
R3252 VSS.n3371 VSS.n3370 185
R3253 VSS.n3373 VSS.n3372 185
R3254 VSS.n3375 VSS.n3374 185
R3255 VSS.n3377 VSS.n3376 185
R3256 VSS.n3379 VSS.n3378 185
R3257 VSS.n3381 VSS.n3380 185
R3258 VSS.n3300 VSS.n1518 185
R3259 VSS.t46 VSS.n1518 185
R3260 VSS.n3299 VSS.n3298 185
R3261 VSS.n3397 VSS.n3396 185
R3262 VSS.n3399 VSS.n3398 185
R3263 VSS.n3290 VSS.n3289 185
R3264 VSS.n3288 VSS.n3287 185
R3265 VSS.n3411 VSS.n3410 185
R3266 VSS.n3413 VSS.n3412 185
R3267 VSS.n3279 VSS.n3278 185
R3268 VSS.n3301 VSS.n3297 185
R3269 VSS.n3389 VSS.n3388 185
R3270 VSS.n3389 VSS.t32 185
R3271 VSS.n3395 VSS.n3394 185
R3272 VSS.n3392 VSS.n3291 185
R3273 VSS.n3391 VSS.n3390 185
R3274 VSS.n3406 VSS.n3405 185
R3275 VSS.n3409 VSS.n3408 185
R3276 VSS.n3280 VSS.n3277 185
R3277 VSS.n3932 VSS.n3931 185
R3278 VSS.n3860 VSS.n1039 185
R3279 VSS.t61 VSS.n1039 185
R3280 VSS.n3858 VSS.n3857 185
R3281 VSS.n3851 VSS.n3850 185
R3282 VSS.n3849 VSS.n3848 185
R3283 VSS.n3842 VSS.n3841 185
R3284 VSS.n3840 VSS.n3839 185
R3285 VSS.n4784 VSS.n4783 185
R3286 VSS.n4786 VSS.n4785 185
R3287 VSS.n1058 VSS.n1057 185
R3288 VSS.n3831 VSS.n3830 185
R3289 VSS.n3859 VSS.n1074 185
R3290 VSS.t50 VSS.n1074 185
R3291 VSS.n3833 VSS.n3832 185
R3292 VSS.n3836 VSS.n3834 185
R3293 VSS.n3838 VSS.n3837 185
R3294 VSS.n3835 VSS.n1066 185
R3295 VSS.n4782 VSS.n4781 185
R3296 VSS.n1067 VSS.n1063 185
R3297 VSS.n1080 VSS.n1062 185
R3298 VSS.n2120 VSS.n2119 185
R3299 VSS.n2118 VSS.n2117 185
R3300 VSS.n2116 VSS.n2115 185
R3301 VSS.n2114 VSS.n2113 185
R3302 VSS.n2112 VSS.n2111 185
R3303 VSS.n2110 VSS.n2109 185
R3304 VSS.n2108 VSS.n2107 185
R3305 VSS.n2106 VSS.n2105 185
R3306 VSS.n2104 VSS.n2045 185
R3307 VSS.n2659 VSS.n2658 185
R3308 VSS.n2661 VSS.n2660 185
R3309 VSS.n2663 VSS.n2662 185
R3310 VSS.n2665 VSS.n2664 185
R3311 VSS.n2667 VSS.n2666 185
R3312 VSS.n2669 VSS.n2668 185
R3313 VSS.n2671 VSS.n2670 185
R3314 VSS.n2673 VSS.n2672 185
R3315 VSS.n2674 VSS.n2063 185
R3316 VSS.n2751 VSS.n2750 185
R3317 VSS.n2750 VSS.t37 185
R3318 VSS.n2044 VSS.n2042 185
R3319 VSS.n2638 VSS.n2637 185
R3320 VSS.n2636 VSS.n2634 185
R3321 VSS.n2646 VSS.n2645 185
R3322 VSS.n2648 VSS.n2647 185
R3323 VSS.n2632 VSS.n2631 185
R3324 VSS.n2630 VSS.n2586 185
R3325 VSS.n2657 VSS.n2656 185
R3326 VSS.n3057 VSS.n3056 185
R3327 VSS.n3056 VSS.t74 185
R3328 VSS.n2001 VSS.n1999 185
R3329 VSS.n2807 VSS.n2806 185
R3330 VSS.n2805 VSS.n2803 185
R3331 VSS.n2815 VSS.n2814 185
R3332 VSS.n2817 VSS.n2816 185
R3333 VSS.n2801 VSS.n2800 185
R3334 VSS.n2799 VSS.n2031 185
R3335 VSS.n2826 VSS.n2825 185
R3336 VSS.n3143 VSS.n1096 185
R3337 VSS.t71 VSS.n1096 185
R3338 VSS.n3141 VSS.n3140 185
R3339 VSS.n3138 VSS.n3137 185
R3340 VSS.n3136 VSS.n3135 185
R3341 VSS.n3124 VSS.n1984 185
R3342 VSS.n3126 VSS.n3125 185
R3343 VSS.n3122 VSS.n3121 185
R3344 VSS.n3120 VSS.n3119 185
R3345 VSS.n3107 VSS.n1990 185
R3346 VSS.n3226 VSS.n1930 185
R3347 VSS.t47 VSS.n1930 185
R3348 VSS.n3229 VSS.n3228 185
R3349 VSS.n3202 VSS.n3201 185
R3350 VSS.n3200 VSS.n3195 185
R3351 VSS.n3238 VSS.n3237 185
R3352 VSS.n3240 VSS.n3239 185
R3353 VSS.n3193 VSS.n3192 185
R3354 VSS.n3191 VSS.n1955 185
R3355 VSS.n3249 VSS.n3248 185
R3356 VSS.n4129 VSS.n1816 185
R3357 VSS.t60 VSS.n1816 185
R3358 VSS.n4127 VSS.n4126 185
R3359 VSS.n4115 VSS.n1902 185
R3360 VSS.n4117 VSS.n4116 185
R3361 VSS.n4113 VSS.n4112 185
R3362 VSS.n4111 VSS.n4110 185
R3363 VSS.n4099 VSS.n1906 185
R3364 VSS.n4101 VSS.n4100 185
R3365 VSS.n4097 VSS.n4096 185
R3366 VSS.n2168 VSS.n2122 185
R3367 VSS.n2166 VSS.n2165 185
R3368 VSS.n2150 VSS.n2123 185
R3369 VSS.n2145 VSS.n2144 185
R3370 VSS.n2142 VSS.n2140 185
R3371 VSS.n2135 VSS.n2071 185
R3372 VSS.n2741 VSS.n2740 185
R3373 VSS.n2738 VSS.n2065 185
R3374 VSS.n2737 VSS.n2064 185
R3375 VSS.n2737 VSS.t57 185
R3376 VSS.n2947 VSS.n2901 185
R3377 VSS.n2945 VSS.n2944 185
R3378 VSS.n2929 VSS.n2902 185
R3379 VSS.n2924 VSS.n2923 185
R3380 VSS.n2921 VSS.n2919 185
R3381 VSS.n2914 VSS.n2028 185
R3382 VSS.n3047 VSS.n3046 185
R3383 VSS.n3044 VSS.n2022 185
R3384 VSS.n3043 VSS.n2021 185
R3385 VSS.n3043 VSS.t52 185
R3386 VSS.n3414 VSS.n1152 185
R3387 VSS.n4743 VSS.n4742 185
R3388 VSS.n4745 VSS.n4744 185
R3389 VSS.n1145 VSS.n1144 185
R3390 VSS.n1143 VSS.n1137 185
R3391 VSS.n4756 VSS.n4755 185
R3392 VSS.n4758 VSS.n4757 185
R3393 VSS.n1092 VSS.n1087 185
R3394 VSS.n4779 VSS.n4778 185
R3395 VSS.t50 VSS.n4779 185
R3396 VSS.n3344 VSS.n1924 185
R3397 VSS.n3342 VSS.n3341 185
R3398 VSS.n3332 VSS.n3306 185
R3399 VSS.n3327 VSS.n3326 185
R3400 VSS.n3324 VSS.n3322 185
R3401 VSS.n3317 VSS.n1952 185
R3402 VSS.n3955 VSS.n3954 185
R3403 VSS.n3952 VSS.n1946 185
R3404 VSS.n3951 VSS.n1945 185
R3405 VSS.n3951 VSS.t32 185
R3406 VSS.n4221 VSS.n1794 185
R3407 VSS.t51 VSS.n1794 185
R3408 VSS.n1846 VSS.n1845 185
R3409 VSS.n4233 VSS.n4232 185
R3410 VSS.n4231 VSS.n4230 185
R3411 VSS.n4245 VSS.n4244 185
R3412 VSS.n4243 VSS.n4242 185
R3413 VSS.n1838 VSS.n1809 185
R3414 VSS.n4280 VSS.n4279 185
R3415 VSS.t51 VSS.n4280 185
R3416 VSS.n1835 VSS.n1808 185
R3417 VSS.n2162 VSS.n2161 185
R3418 VSS.n2164 VSS.n2163 185
R3419 VSS.n2149 VSS.n2148 185
R3420 VSS.n2147 VSS.n2146 185
R3421 VSS.n2139 VSS.n2138 185
R3422 VSS.n2137 VSS.n2136 185
R3423 VSS.n2070 VSS.n2069 185
R3424 VSS.n2068 VSS.n2046 185
R3425 VSS.t37 VSS.n2046 185
R3426 VSS.n2748 VSS.n2747 185
R3427 VSS.n2941 VSS.n2940 185
R3428 VSS.n2943 VSS.n2942 185
R3429 VSS.n2928 VSS.n2927 185
R3430 VSS.n2926 VSS.n2925 185
R3431 VSS.n2918 VSS.n2917 185
R3432 VSS.n2916 VSS.n2915 185
R3433 VSS.n2027 VSS.n2026 185
R3434 VSS.n2025 VSS.n2003 185
R3435 VSS.t74 VSS.n2003 185
R3436 VSS.n3054 VSS.n3053 185
R3437 VSS.n4739 VSS.n4738 185
R3438 VSS.n4741 VSS.n4740 185
R3439 VSS.n1149 VSS.n1148 185
R3440 VSS.n1147 VSS.n1146 185
R3441 VSS.n4752 VSS.n4751 185
R3442 VSS.n4754 VSS.n4753 185
R3443 VSS.n1134 VSS.n1091 185
R3444 VSS.n4775 VSS.n1093 185
R3445 VSS.n4775 VSS.t71 185
R3446 VSS.n4777 VSS.n4776 185
R3447 VSS.n3966 VSS.n3965 185
R3448 VSS.n3340 VSS.n1925 185
R3449 VSS.n3331 VSS.n3330 185
R3450 VSS.n3329 VSS.n3328 185
R3451 VSS.n3321 VSS.n3320 185
R3452 VSS.n3319 VSS.n3318 185
R3453 VSS.n1951 VSS.n1950 185
R3454 VSS.n1949 VSS.n1927 185
R3455 VSS.t47 VSS.n1927 185
R3456 VSS.n3962 VSS.n3961 185
R3457 VSS.n4220 VSS.n4219 185
R3458 VSS.n4218 VSS.n1848 185
R3459 VSS.n4229 VSS.n4228 185
R3460 VSS.n4227 VSS.n1844 185
R3461 VSS.n4241 VSS.n4240 185
R3462 VSS.n4239 VSS.n1842 185
R3463 VSS.n1839 VSS.n1813 185
R3464 VSS.n4278 VSS.n4277 185
R3465 VSS.n4277 VSS.t60 185
R3466 VSS.n1834 VSS.n1812 185
R3467 VSS.n4272 VSS.n4271 185
R3468 VSS.n4270 VSS.n4269 185
R3469 VSS.n4268 VSS.n4267 185
R3470 VSS.n4266 VSS.n4265 185
R3471 VSS.n4264 VSS.n4263 185
R3472 VSS.n4262 VSS.n4261 185
R3473 VSS.n4260 VSS.n4259 185
R3474 VSS.n4258 VSS.n4257 185
R3475 VSS.n4281 VSS.n1779 185
R3476 VSS.n4297 VSS.n1777 185
R3477 VSS.n4336 VSS.n4335 185
R3478 VSS.n4334 VSS.n1778 185
R3479 VSS.n4333 VSS.n4332 185
R3480 VSS.n4331 VSS.n4330 185
R3481 VSS.n4329 VSS.n4328 185
R3482 VSS.n4327 VSS.n4326 185
R3483 VSS.n4325 VSS.n4324 185
R3484 VSS.n4323 VSS.n4322 185
R3485 VSS.n2479 VSS.n2453 185
R3486 VSS.n2481 VSS.n2480 185
R3487 VSS.n2473 VSS.n2472 185
R3488 VSS.n2471 VSS.n2470 185
R3489 VSS.n2464 VSS.n2463 185
R3490 VSS.n2462 VSS.n2461 185
R3491 VSS.n4288 VSS.n4287 185
R3492 VSS.n4290 VSS.n4289 185
R3493 VSS.n1782 VSS.n1781 185
R3494 VSS.n2488 VSS.n2487 185
R3495 VSS.n2486 VSS.n2485 185
R3496 VSS.n2455 VSS.n2454 185
R3497 VSS.n2457 VSS.n2456 185
R3498 VSS.n2460 VSS.n2459 185
R3499 VSS.n2458 VSS.n1791 185
R3500 VSS.n4286 VSS.n4285 185
R3501 VSS.n1790 VSS.n1784 185
R3502 VSS.n4282 VSS.n1783 185
R3503 VSS.n2508 VSS.n2507 185
R3504 VSS.n2506 VSS.n2505 185
R3505 VSS.n2504 VSS.n2503 185
R3506 VSS.n2502 VSS.n2501 185
R3507 VSS.n2500 VSS.n2499 185
R3508 VSS.n2498 VSS.n2497 185
R3509 VSS.n2496 VSS.n2495 185
R3510 VSS.n2494 VSS.n2493 185
R3511 VSS.n2492 VSS.n2491 185
R3512 VSS.n1739 VSS.n1408 185
R3513 VSS.n2394 VSS.n2393 185
R3514 VSS.n2396 VSS.n2395 185
R3515 VSS.n2398 VSS.n2397 185
R3516 VSS.n2400 VSS.n2399 185
R3517 VSS.n2402 VSS.n2401 185
R3518 VSS.n2404 VSS.n2403 185
R3519 VSS.n2406 VSS.n2405 185
R3520 VSS.n2408 VSS.n2407 185
R3521 VSS.n532 VSS.n290 185
R3522 VSS.n5264 VSS.n5263 185
R3523 VSS.n5266 VSS.n5265 185
R3524 VSS.n283 VSS.n282 185
R3525 VSS.n281 VSS.n275 185
R3526 VSS.n5277 VSS.n5276 185
R3527 VSS.n5279 VSS.n5278 185
R3528 VSS.n245 VSS.n240 185
R3529 VSS.n5310 VSS.n5309 185
R3530 VSS.t39 VSS.n5310 185
R3531 VSS.n891 VSS.n718 185
R3532 VSS.n5057 VSS.n5056 185
R3533 VSS.n5059 VSS.n5058 185
R3534 VSS.n711 VSS.n710 185
R3535 VSS.n709 VSS.n703 185
R3536 VSS.n5070 VSS.n5069 185
R3537 VSS.n5072 VSS.n5071 185
R3538 VSS.n494 VSS.n489 185
R3539 VSS.n5103 VSS.n5102 185
R3540 VSS.t73 VSS.n5103 185
R3541 VSS.n3804 VSS.n3803 185
R3542 VSS.n3798 VSS.n3797 185
R3543 VSS.n3796 VSS.n3795 185
R3544 VSS.n3790 VSS.n3789 185
R3545 VSS.n3788 VSS.n3787 185
R3546 VSS.n3782 VSS.n3781 185
R3547 VSS.n3780 VSS.n3779 185
R3548 VSS.n1035 VSS.n1030 185
R3549 VSS.n4850 VSS.n4849 185
R3550 VSS.t69 VSS.n4850 185
R3551 VSS.n1585 VSS.n1555 185
R3552 VSS.n4431 VSS.n4430 185
R3553 VSS.n4433 VSS.n4432 185
R3554 VSS.n1548 VSS.n1547 185
R3555 VSS.n1546 VSS.n1540 185
R3556 VSS.n4444 VSS.n4443 185
R3557 VSS.n4446 VSS.n4445 185
R3558 VSS.n1514 VSS.n1509 185
R3559 VSS.n4477 VSS.n4476 185
R3560 VSS.t49 VSS.n4477 185
R3561 VSS.n2434 VSS.n2433 185
R3562 VSS.n2432 VSS.n2431 185
R3563 VSS.n2426 VSS.n2425 185
R3564 VSS.n2424 VSS.n2423 185
R3565 VSS.n4347 VSS.n4346 185
R3566 VSS.n4345 VSS.n4344 185
R3567 VSS.n1757 VSS.n1756 185
R3568 VSS.n1755 VSS.n1749 185
R3569 VSS.n4360 VSS.n4359 185
R3570 VSS.n5260 VSS.n5259 185
R3571 VSS.n5262 VSS.n5261 185
R3572 VSS.n287 VSS.n286 185
R3573 VSS.n285 VSS.n284 185
R3574 VSS.n5273 VSS.n5272 185
R3575 VSS.n5275 VSS.n5274 185
R3576 VSS.n272 VSS.n244 185
R3577 VSS.n5306 VSS.n246 185
R3578 VSS.n5306 VSS.t30 185
R3579 VSS.n5308 VSS.n5307 185
R3580 VSS.n5053 VSS.n5052 185
R3581 VSS.n5055 VSS.n5054 185
R3582 VSS.n715 VSS.n714 185
R3583 VSS.n713 VSS.n712 185
R3584 VSS.n5066 VSS.n5065 185
R3585 VSS.n5068 VSS.n5067 185
R3586 VSS.n700 VSS.n493 185
R3587 VSS.n5099 VSS.n495 185
R3588 VSS.n5099 VSS.t59 185
R3589 VSS.n5101 VSS.n5100 185
R3590 VSS.n3799 VSS.n3754 185
R3591 VSS.n3801 VSS.n3800 185
R3592 VSS.n3794 VSS.n3793 185
R3593 VSS.n3792 VSS.n3791 185
R3594 VSS.n3786 VSS.n3785 185
R3595 VSS.n3784 VSS.n3783 185
R3596 VSS.n3778 VSS.n1034 185
R3597 VSS.n4846 VSS.n1036 185
R3598 VSS.n4846 VSS.t61 185
R3599 VSS.n4848 VSS.n4847 185
R3600 VSS.n4427 VSS.n4426 185
R3601 VSS.n4429 VSS.n4428 185
R3602 VSS.n1552 VSS.n1551 185
R3603 VSS.n1550 VSS.n1549 185
R3604 VSS.n4440 VSS.n4439 185
R3605 VSS.n4442 VSS.n4441 185
R3606 VSS.n1537 VSS.n1513 185
R3607 VSS.n4473 VSS.n1515 185
R3608 VSS.n4473 VSS.t46 185
R3609 VSS.n4475 VSS.n4474 185
R3610 VSS.n2510 VSS.n2509 185
R3611 VSS.n2430 VSS.n2429 185
R3612 VSS.n2428 VSS.n2427 185
R3613 VSS.n2422 VSS.n1762 185
R3614 VSS.n4343 VSS.n4342 185
R3615 VSS.n4340 VSS.n1761 185
R3616 VSS.n4339 VSS.n4338 185
R3617 VSS.n4356 VSS.n4355 185
R3618 VSS.n4358 VSS.n4357 185
R3619 VSS.n5417 VSS.n5416 185
R3620 VSS.n5393 VSS.n103 185
R3621 VSS.n5392 VSS.n5391 185
R3622 VSS.n5390 VSS.n5389 185
R3623 VSS.n5402 VSS.n5401 185
R3624 VSS.n5404 VSS.n5403 185
R3625 VSS.n132 VSS.n131 185
R3626 VSS.n124 VSS.n105 185
R3627 VSS.t41 VSS.n105 185
R3628 VSS.n5413 VSS.n5412 185
R3629 VSS.n5204 VSS.n5203 185
R3630 VSS.n5180 VSS.n402 185
R3631 VSS.n5179 VSS.n5178 185
R3632 VSS.n5177 VSS.n5176 185
R3633 VSS.n5189 VSS.n5188 185
R3634 VSS.n5191 VSS.n5190 185
R3635 VSS.n5170 VSS.n5169 185
R3636 VSS.n5160 VSS.n404 185
R3637 VSS.t53 VSS.n404 185
R3638 VSS.n5200 VSS.n5199 185
R3639 VSS.n4951 VSS.n4950 185
R3640 VSS.n4927 VSS.n817 185
R3641 VSS.n4926 VSS.n4925 185
R3642 VSS.n4924 VSS.n4923 185
R3643 VSS.n4936 VSS.n4935 185
R3644 VSS.n4938 VSS.n4937 185
R3645 VSS.n4917 VSS.n4916 185
R3646 VSS.n4907 VSS.n819 185
R3647 VSS.t65 VSS.n819 185
R3648 VSS.n4947 VSS.n4946 185
R3649 VSS.n3647 VSS.n3646 185
R3650 VSS.n3649 VSS.n3648 185
R3651 VSS.n3643 VSS.n3642 185
R3652 VSS.n3641 VSS.n3640 185
R3653 VSS.n3658 VSS.n3657 185
R3654 VSS.n3660 VSS.n3659 185
R3655 VSS.n3634 VSS.n3633 185
R3656 VSS.n3624 VSS.n3488 185
R3657 VSS.t54 VSS.n3488 185
R3658 VSS.n3669 VSS.n3668 185
R3659 VSS.n43 VSS.n36 185
R3660 VSS.n5505 VSS.n5504 185
R3661 VSS.n5502 VSS.n40 185
R3662 VSS.n5501 VSS.n45 185
R3663 VSS.n5499 VSS.n5498 185
R3664 VSS.n49 VSS.n46 185
R3665 VSS.n5486 VSS.n5485 185
R3666 VSS.n5488 VSS.n5487 185
R3667 VSS.n5487 VSS.t56 185
R3668 VSS.n5483 VSS.n53 185
R3669 VSS.n5538 VSS.n19 175.546
R3670 VSS.n5542 VSS.n19 175.546
R3671 VSS.n5542 VSS.n17 175.546
R3672 VSS.n5546 VSS.n17 175.546
R3673 VSS.n5546 VSS.n12 175.546
R3674 VSS.n5550 VSS.n12 175.546
R3675 VSS.n5550 VSS.n10 175.546
R3676 VSS.n5555 VSS.n10 175.546
R3677 VSS.n5555 VSS.n7 175.546
R3678 VSS.n5559 VSS.n7 175.546
R3679 VSS.n5560 VSS.n5559 175.546
R3680 VSS.n4587 VSS.n1388 175.546
R3681 VSS.n4587 VSS.n1405 175.546
R3682 VSS.n4615 VSS.n1405 175.546
R3683 VSS.n4615 VSS.n1406 175.546
R3684 VSS.n4611 VSS.n1406 175.546
R3685 VSS.n4611 VSS.n4609 175.546
R3686 VSS.n4609 VSS.n4591 175.546
R3687 VSS.n4605 VSS.n4591 175.546
R3688 VSS.n4605 VSS.n4593 175.546
R3689 VSS.n4601 VSS.n4593 175.546
R3690 VSS.n4601 VSS.n4597 175.546
R3691 VSS.n2541 VSS.n2540 175.546
R3692 VSS.n2540 VSS.n2517 175.546
R3693 VSS.n2536 VSS.n2517 175.546
R3694 VSS.n2536 VSS.n1380 175.546
R3695 VSS.n4655 VSS.n1380 175.546
R3696 VSS.n4655 VSS.n1381 175.546
R3697 VSS.n4651 VSS.n1381 175.546
R3698 VSS.n4651 VSS.n1384 175.546
R3699 VSS.n4647 VSS.n1384 175.546
R3700 VSS.n4647 VSS.n1386 175.546
R3701 VSS.n4678 VSS.n1362 175.546
R3702 VSS.n4674 VSS.n1362 175.546
R3703 VSS.n4674 VSS.n1364 175.546
R3704 VSS.n4670 VSS.n1364 175.546
R3705 VSS.n4670 VSS.n4667 175.546
R3706 VSS.n4667 VSS.n4666 175.546
R3707 VSS.n4666 VSS.n1366 175.546
R3708 VSS.n2524 VSS.n1366 175.546
R3709 VSS.n2524 VSS.n2519 175.546
R3710 VSS.n2529 VSS.n2519 175.546
R3711 VSS.n2529 VSS.n2521 175.546
R3712 VSS.n4209 VSS.n1855 175.546
R3713 VSS.n4209 VSS.n1856 175.546
R3714 VSS.n4205 VSS.n1856 175.546
R3715 VSS.n4205 VSS.n4184 175.546
R3716 VSS.n4201 VSS.n4184 175.546
R3717 VSS.n4201 VSS.n4200 175.546
R3718 VSS.n4200 VSS.n4186 175.546
R3719 VSS.n4196 VSS.n4186 175.546
R3720 VSS.n4196 VSS.n4188 175.546
R3721 VSS.n4192 VSS.n4188 175.546
R3722 VSS.n2321 VSS.n2268 175.546
R3723 VSS.n2321 VSS.n2269 175.546
R3724 VSS.n2317 VSS.n2269 175.546
R3725 VSS.n2317 VSS.n2272 175.546
R3726 VSS.n2313 VSS.n2272 175.546
R3727 VSS.n2313 VSS.n2274 175.546
R3728 VSS.n2309 VSS.n2274 175.546
R3729 VSS.n2309 VSS.n2276 175.546
R3730 VSS.n2305 VSS.n2276 175.546
R3731 VSS.n2305 VSS.n2278 175.546
R3732 VSS.n2386 VSS.n2385 175.546
R3733 VSS.n2385 VSS.n2255 175.546
R3734 VSS.n2381 VSS.n2255 175.546
R3735 VSS.n2381 VSS.n2258 175.546
R3736 VSS.n2377 VSS.n2258 175.546
R3737 VSS.n2377 VSS.n2261 175.546
R3738 VSS.n2373 VSS.n2261 175.546
R3739 VSS.n2373 VSS.n2263 175.546
R3740 VSS.n2369 VSS.n2263 175.546
R3741 VSS.n2369 VSS.n2366 175.546
R3742 VSS.n2570 VSS.n2241 175.546
R3743 VSS.n2566 VSS.n2241 175.546
R3744 VSS.n2566 VSS.n2243 175.546
R3745 VSS.n2562 VSS.n2243 175.546
R3746 VSS.n2562 VSS.n2559 175.546
R3747 VSS.n2559 VSS.n2558 175.546
R3748 VSS.n2558 VSS.n2246 175.546
R3749 VSS.n2554 VSS.n2246 175.546
R3750 VSS.n2554 VSS.n2249 175.546
R3751 VSS.n2550 VSS.n2249 175.546
R3752 VSS.n2550 VSS.n2253 175.546
R3753 VSS.n2686 VSS.n2580 175.546
R3754 VSS.n2686 VSS.n2578 175.546
R3755 VSS.n2690 VSS.n2578 175.546
R3756 VSS.n2690 VSS.n2576 175.546
R3757 VSS.n2694 VSS.n2576 175.546
R3758 VSS.n2695 VSS.n2694 175.546
R3759 VSS.n2698 VSS.n2695 175.546
R3760 VSS.n2698 VSS.n2574 175.546
R3761 VSS.n2703 VSS.n2574 175.546
R3762 VSS.n2703 VSS.n2571 175.546
R3763 VSS.n2296 VSS.n2285 175.546
R3764 VSS.n2292 VSS.n2285 175.546
R3765 VSS.n2292 VSS.n2288 175.546
R3766 VSS.n2288 VSS.n160 175.546
R3767 VSS.n5384 VSS.n160 175.546
R3768 VSS.n5384 VSS.n161 175.546
R3769 VSS.n5380 VSS.n161 175.546
R3770 VSS.n5380 VSS.n164 175.546
R3771 VSS.n5376 VSS.n164 175.546
R3772 VSS.n5376 VSS.n166 175.546
R3773 VSS.n2620 VSS.n2592 175.546
R3774 VSS.n2616 VSS.n2592 175.546
R3775 VSS.n2616 VSS.n2594 175.546
R3776 VSS.n2612 VSS.n2594 175.546
R3777 VSS.n2612 VSS.n2610 175.546
R3778 VSS.n2610 VSS.n2596 175.546
R3779 VSS.n2606 VSS.n2596 175.546
R3780 VSS.n2606 VSS.n2602 175.546
R3781 VSS.n2602 VSS.n2601 175.546
R3782 VSS.n2601 VSS.n2598 175.546
R3783 VSS.n2624 VSS.n2587 175.546
R3784 VSS.n2654 VSS.n2587 175.546
R3785 VSS.n2654 VSS.n2588 175.546
R3786 VSS.n2650 VSS.n2588 175.546
R3787 VSS.n2650 VSS.n2628 175.546
R3788 VSS.n2643 VSS.n2628 175.546
R3789 VSS.n2643 VSS.n2640 175.546
R3790 VSS.n2640 VSS.n2041 175.546
R3791 VSS.n2753 VSS.n2041 175.546
R3792 VSS.n2753 VSS.n2039 175.546
R3793 VSS.n2757 VSS.n2039 175.546
R3794 VSS.n5372 VSS.n125 175.546
R3795 VSS.n5410 VSS.n125 175.546
R3796 VSS.n5410 VSS.n126 175.546
R3797 VSS.n5406 VSS.n126 175.546
R3798 VSS.n5406 VSS.n129 175.546
R3799 VSS.n5399 VSS.n129 175.546
R3800 VSS.n5399 VSS.n134 175.546
R3801 VSS.n5395 VSS.n134 175.546
R3802 VSS.n5395 VSS.n5387 175.546
R3803 VSS.n5387 VSS.n100 175.546
R3804 VSS.n5422 VSS.n100 175.546
R3805 VSS.n5476 VSS.n52 175.546
R3806 VSS.n5490 VSS.n52 175.546
R3807 VSS.n5490 VSS.n48 175.546
R3808 VSS.n5494 VSS.n48 175.546
R3809 VSS.n5495 VSS.n5494 175.546
R3810 VSS.n5496 VSS.n5495 175.546
R3811 VSS.n5496 VSS.n39 175.546
R3812 VSS.n5507 VSS.n39 175.546
R3813 VSS.n5507 VSS.n37 175.546
R3814 VSS.n5511 VSS.n37 175.546
R3815 VSS.n5511 VSS.n5 175.546
R3816 VSS.n5163 VSS.n5161 175.546
R3817 VSS.n5197 VSS.n5161 175.546
R3818 VSS.n5197 VSS.n5162 175.546
R3819 VSS.n5193 VSS.n5162 175.546
R3820 VSS.n5193 VSS.n5167 175.546
R3821 VSS.n5186 VSS.n5167 175.546
R3822 VSS.n5186 VSS.n5172 175.546
R3823 VSS.n5182 VSS.n5172 175.546
R3824 VSS.n5182 VSS.n5174 175.546
R3825 VSS.n5174 VSS.n399 175.546
R3826 VSS.n5209 VSS.n399 175.546
R3827 VSS.n3627 VSS.n3625 175.546
R3828 VSS.n3666 VSS.n3625 175.546
R3829 VSS.n3666 VSS.n3626 175.546
R3830 VSS.n3662 VSS.n3626 175.546
R3831 VSS.n3662 VSS.n3631 175.546
R3832 VSS.n3655 VSS.n3631 175.546
R3833 VSS.n3655 VSS.n3636 175.546
R3834 VSS.n3651 VSS.n3636 175.546
R3835 VSS.n3651 VSS.n3638 175.546
R3836 VSS.n3638 VSS.n61 175.546
R3837 VSS.n5470 VSS.n61 175.546
R3838 VSS.n4910 VSS.n4908 175.546
R3839 VSS.n4944 VSS.n4908 175.546
R3840 VSS.n4944 VSS.n4909 175.546
R3841 VSS.n4940 VSS.n4909 175.546
R3842 VSS.n4940 VSS.n4914 175.546
R3843 VSS.n4933 VSS.n4914 175.546
R3844 VSS.n4933 VSS.n4919 175.546
R3845 VSS.n4929 VSS.n4919 175.546
R3846 VSS.n4929 VSS.n4921 175.546
R3847 VSS.n4921 VSS.n814 175.546
R3848 VSS.n4956 VSS.n814 175.546
R3849 VSS.n2793 VSS.n2032 175.546
R3850 VSS.n2823 VSS.n2032 175.546
R3851 VSS.n2823 VSS.n2033 175.546
R3852 VSS.n2819 VSS.n2033 175.546
R3853 VSS.n2819 VSS.n2797 175.546
R3854 VSS.n2812 VSS.n2797 175.546
R3855 VSS.n2812 VSS.n2809 175.546
R3856 VSS.n2809 VSS.n1998 175.546
R3857 VSS.n3059 VSS.n1998 175.546
R3858 VSS.n3059 VSS.n1996 175.546
R3859 VSS.n3063 VSS.n1996 175.546
R3860 VSS.n3113 VSS.n1991 175.546
R3861 VSS.n3117 VSS.n1991 175.546
R3862 VSS.n3117 VSS.n1988 175.546
R3863 VSS.n3128 VSS.n1988 175.546
R3864 VSS.n3128 VSS.n1985 175.546
R3865 VSS.n3133 VSS.n1985 175.546
R3866 VSS.n3133 VSS.n1986 175.546
R3867 VSS.n1986 VSS.n1982 175.546
R3868 VSS.n3145 VSS.n1982 175.546
R3869 VSS.n3145 VSS.n1980 175.546
R3870 VSS.n3149 VSS.n1980 175.546
R3871 VSS.n4157 VSS.n1867 175.546
R3872 VSS.n4162 VSS.n1867 175.546
R3873 VSS.n4162 VSS.n1865 175.546
R3874 VSS.n4166 VSS.n1865 175.546
R3875 VSS.n4166 VSS.n1863 175.546
R3876 VSS.n4171 VSS.n1863 175.546
R3877 VSS.n4171 VSS.n1860 175.546
R3878 VSS.n4175 VSS.n1860 175.546
R3879 VSS.n4176 VSS.n4175 175.546
R3880 VSS.n4177 VSS.n4176 175.546
R3881 VSS.n4079 VSS.n1909 175.546
R3882 VSS.n4103 VSS.n1909 175.546
R3883 VSS.n4103 VSS.n1907 175.546
R3884 VSS.n4108 VSS.n1907 175.546
R3885 VSS.n4108 VSS.n1904 175.546
R3886 VSS.n4119 VSS.n1904 175.546
R3887 VSS.n4119 VSS.n1903 175.546
R3888 VSS.n4124 VSS.n1903 175.546
R3889 VSS.n4124 VSS.n1901 175.546
R3890 VSS.n4150 VSS.n1901 175.546
R3891 VSS.n4151 VSS.n4150 175.546
R3892 VSS.n3185 VSS.n1956 175.546
R3893 VSS.n3246 VSS.n1956 175.546
R3894 VSS.n3246 VSS.n1957 175.546
R3895 VSS.n3242 VSS.n1957 175.546
R3896 VSS.n3242 VSS.n3189 175.546
R3897 VSS.n3235 VSS.n3189 175.546
R3898 VSS.n3235 VSS.n3196 175.546
R3899 VSS.n3231 VSS.n3196 175.546
R3900 VSS.n3231 VSS.n3198 175.546
R3901 VSS.n3224 VSS.n3198 175.546
R3902 VSS.n3224 VSS.n1912 175.546
R3903 VSS.n4664 VSS.n1368 167.089
R3904 VSS.n4640 VSS.t6 167.089
R3905 VSS.n2509 VSS.n2508 163.333
R3906 VSS.n959 VSS.n958 163.333
R3907 VSS.n1434 VSS.n1433 163.333
R3908 VSS.n1739 VSS.n1738 163.333
R3909 VSS.n4499 VSS.n4498 163.333
R3910 VSS.n3687 VSS.n3686 163.333
R3911 VSS.n1881 VSS.n1874 161.972
R3912 VSS.n1358 VSS.n1265 160.662
R3913 VSS.n2545 VSS.n2390 160.662
R3914 VSS.n4642 VSS.n4641 160.662
R3915 VSS.n4598 VSS.n20 160.662
R3916 VSS.n4289 VSS.n4288 150
R3917 VSS.n2463 VSS.n2462 150
R3918 VSS.n2472 VSS.n2471 150
R3919 VSS.n2480 VSS.n2479 150
R3920 VSS.n2493 VSS.n2492 150
R3921 VSS.n2497 VSS.n2496 150
R3922 VSS.n2501 VSS.n2500 150
R3923 VSS.n2505 VSS.n2504 150
R3924 VSS.n4357 VSS.n4356 150
R3925 VSS.n4340 VSS.n4339 150
R3926 VSS.n4342 VSS.n1762 150
R3927 VSS.n2429 VSS.n2428 150
R3928 VSS.n4336 VSS.n1778 150
R3929 VSS.n4332 VSS.n4331 150
R3930 VSS.n4328 VSS.n4327 150
R3931 VSS.n4324 VSS.n4323 150
R3932 VSS.n4280 VSS.n1808 150
R3933 VSS.n4280 VSS.n1809 150
R3934 VSS.n4244 VSS.n4243 150
R3935 VSS.n4232 VSS.n4231 150
R3936 VSS.n1845 VSS.n1794 150
R3937 VSS.n4271 VSS.n4270 150
R3938 VSS.n4267 VSS.n4266 150
R3939 VSS.n4263 VSS.n4262 150
R3940 VSS.n4259 VSS.n4258 150
R3941 VSS.n4285 VSS.n1790 150
R3942 VSS.n2459 VSS.n1791 150
R3943 VSS.n2456 VSS.n2455 150
R3944 VSS.n2487 VSS.n2486 150
R3945 VSS.n2439 VSS.n2438 150
R3946 VSS.n2443 VSS.n2442 150
R3947 VSS.n2447 VSS.n2446 150
R3948 VSS.n2451 VSS.n2450 150
R3949 VSS.n4100 VSS.n4099 150
R3950 VSS.n4112 VSS.n4111 150
R3951 VSS.n4116 VSS.n4115 150
R3952 VSS.n4126 VSS.n1816 150
R3953 VSS.n4144 VSS.n4143 150
R3954 VSS.n4140 VSS.n4139 150
R3955 VSS.n4136 VSS.n4135 150
R3956 VSS.n4132 VSS.n4131 150
R3957 VSS.n4277 VSS.n1812 150
R3958 VSS.n4277 VSS.n1813 150
R3959 VSS.n4240 VSS.n4239 150
R3960 VSS.n4228 VSS.n4227 150
R3961 VSS.n4219 VSS.n4218 150
R3962 VSS.n4092 VSS.n4091 150
R3963 VSS.n4088 VSS.n4087 150
R3964 VSS.n4084 VSS.n4083 150
R3965 VSS.n4275 VSS.n1831 150
R3966 VSS.n3192 VSS.n3191 150
R3967 VSS.n3239 VSS.n3238 150
R3968 VSS.n3201 VSS.n3200 150
R3969 VSS.n3228 VSS.n1930 150
R3970 VSS.n3216 VSS.n3215 150
R3971 VSS.n3212 VSS.n3211 150
R3972 VSS.n3208 VSS.n3207 150
R3973 VSS.n3204 VSS.n1926 150
R3974 VSS.n3962 VSS.n1927 150
R3975 VSS.n1950 VSS.n1927 150
R3976 VSS.n3320 VSS.n3319 150
R3977 VSS.n3330 VSS.n3329 150
R3978 VSS.n3965 VSS.n1925 150
R3979 VSS.n3254 VSS.n3253 150
R3980 VSS.n3258 VSS.n3257 150
R3981 VSS.n3262 VSS.n3261 150
R3982 VSS.n3264 VSS.n1944 150
R3983 VSS.n3121 VSS.n3120 150
R3984 VSS.n3125 VSS.n3124 150
R3985 VSS.n3137 VSS.n3136 150
R3986 VSS.n3140 VSS.n1096 150
R3987 VSS.n1975 VSS.n1974 150
R3988 VSS.n1971 VSS.n1970 150
R3989 VSS.n1967 VSS.n1966 150
R3990 VSS.n1963 VSS.n1962 150
R3991 VSS.n4776 VSS.n4775 150
R3992 VSS.n4775 VSS.n1091 150
R3993 VSS.n4753 VSS.n4752 150
R3994 VSS.n1148 VSS.n1147 150
R3995 VSS.n4740 VSS.n4739 150
R3996 VSS.n3105 VSS.n3104 150
R3997 VSS.n3101 VSS.n3100 150
R3998 VSS.n4773 VSS.n1111 150
R3999 VSS.n4769 VSS.n1110 150
R4000 VSS.n2800 VSS.n2799 150
R4001 VSS.n2816 VSS.n2815 150
R4002 VSS.n2806 VSS.n2805 150
R4003 VSS.n3056 VSS.n2001 150
R4004 VSS.n2886 VSS.n2885 150
R4005 VSS.n2890 VSS.n2889 150
R4006 VSS.n2894 VSS.n2893 150
R4007 VSS.n2898 VSS.n2897 150
R4008 VSS.n3054 VSS.n2003 150
R4009 VSS.n2026 VSS.n2003 150
R4010 VSS.n2917 VSS.n2916 150
R4011 VSS.n2927 VSS.n2926 150
R4012 VSS.n2942 VSS.n2941 150
R4013 VSS.n2831 VSS.n2830 150
R4014 VSS.n2835 VSS.n2834 150
R4015 VSS.n2839 VSS.n2838 150
R4016 VSS.n2841 VSS.n2020 150
R4017 VSS.n4785 VSS.n4784 150
R4018 VSS.n3841 VSS.n3840 150
R4019 VSS.n3850 VSS.n3849 150
R4020 VSS.n3857 VSS.n1039 150
R4021 VSS.n4844 VSS.n1054 150
R4022 VSS.n4840 VSS.n4839 150
R4023 VSS.n4836 VSS.n4835 150
R4024 VSS.n4832 VSS.n4831 150
R4025 VSS.n4847 VSS.n4846 150
R4026 VSS.n4846 VSS.n1034 150
R4027 VSS.n3785 VSS.n3784 150
R4028 VSS.n3793 VSS.n3792 150
R4029 VSS.n3800 VSS.n3799 150
R4030 VSS.n3826 VSS.n3825 150
R4031 VSS.n3822 VSS.n3821 150
R4032 VSS.n3818 VSS.n3817 150
R4033 VSS.n3814 VSS.n3813 150
R4034 VSS.n4779 VSS.n1087 150
R4035 VSS.n4757 VSS.n4756 150
R4036 VSS.n1144 VSS.n1143 150
R4037 VSS.n4744 VSS.n4743 150
R4038 VSS.n1126 VSS.n1125 150
R4039 VSS.n1122 VSS.n1121 150
R4040 VSS.n1118 VSS.n1117 150
R4041 VSS.n1114 VSS.n1113 150
R4042 VSS.n1080 VSS.n1067 150
R4043 VSS.n4781 VSS.n1066 150
R4044 VSS.n3837 VSS.n3836 150
R4045 VSS.n3832 VSS.n1074 150
R4046 VSS.n3830 VSS.n1074 150
R4047 VSS.n3419 VSS.n3418 150
R4048 VSS.n3423 VSS.n3422 150
R4049 VSS.n3427 VSS.n3426 150
R4050 VSS.n3431 VSS.n3430 150
R4051 VSS.n5310 VSS.n240 150
R4052 VSS.n5278 VSS.n5277 150
R4053 VSS.n282 VSS.n281 150
R4054 VSS.n5265 VSS.n5264 150
R4055 VSS.n2342 VSS.n2341 150
R4056 VSS.n2346 VSS.n2345 150
R4057 VSS.n2350 VSS.n2349 150
R4058 VSS.n2354 VSS.n2353 150
R4059 VSS.n5327 VSS.n5326 150
R4060 VSS.n225 VSS.n224 150
R4061 VSS.n5312 VSS.n219 150
R4062 VSS.n229 VSS.n220 150
R4063 VSS.n613 VSS.n229 150
R4064 VSS.n537 VSS.n536 150
R4065 VSS.n541 VSS.n540 150
R4066 VSS.n545 VSS.n544 150
R4067 VSS.n549 VSS.n548 150
R4068 VSS.n175 VSS.n174 150
R4069 VSS.n5336 VSS.n5335 150
R4070 VSS.n578 VSS.n577 150
R4071 VSS.n585 VSS.n108 150
R4072 VSS.n5355 VSS.n5354 150
R4073 VSS.n5359 VSS.n5358 150
R4074 VSS.n5363 VSS.n5362 150
R4075 VSS.n5365 VSS.n122 150
R4076 VSS.n5413 VSS.n105 150
R4077 VSS.n131 VSS.n105 150
R4078 VSS.n5403 VSS.n5402 150
R4079 VSS.n5391 VSS.n5390 150
R4080 VSS.n5416 VSS.n103 150
R4081 VSS.n563 VSS.n562 150
R4082 VSS.n559 VSS.n558 150
R4083 VSS.n555 VSS.n554 150
R4084 VSS.n551 VSS.n104 150
R4085 VSS.n5330 VSS.n201 150
R4086 VSS.n214 VSS.n213 150
R4087 VSS.n5316 VSS.n5315 150
R4088 VSS.n626 VSS.n625 150
R4089 VSS.n2337 VSS.n2336 150
R4090 VSS.n2333 VSS.n2332 150
R4091 VSS.n2329 VSS.n2328 150
R4092 VSS.n2325 VSS.n2324 150
R4093 VSS.n5347 VSS.n5346 150
R4094 VSS.n184 VSS.n183 150
R4095 VSS.n5332 VSS.n181 150
R4096 VSS.n570 VSS.n190 150
R4097 VSS.n567 VSS.n190 150
R4098 VSS.n610 VSS.n609 150
R4099 VSS.n606 VSS.n605 150
R4100 VSS.n602 VSS.n601 150
R4101 VSS.n598 VSS.n597 150
R4102 VSS.n429 VSS.n428 150
R4103 VSS.n5128 VSS.n5127 150
R4104 VSS.n861 VSS.n860 150
R4105 VSS.n866 VSS.n407 150
R4106 VSS.n887 VSS.n886 150
R4107 VSS.n883 VSS.n882 150
R4108 VSS.n879 VSS.n878 150
R4109 VSS.n875 VSS.n403 150
R4110 VSS.n5200 VSS.n404 150
R4111 VSS.n5169 VSS.n404 150
R4112 VSS.n5190 VSS.n5189 150
R4113 VSS.n5178 VSS.n5177 150
R4114 VSS.n5203 VSS.n402 150
R4115 VSS.n5145 VSS.n5144 150
R4116 VSS.n5149 VSS.n5148 150
R4117 VSS.n5153 VSS.n5152 150
R4118 VSS.n5155 VSS.n421 150
R4119 VSS.n463 VSS.n456 150
R4120 VSS.n5109 VSS.n5108 150
R4121 VSS.n924 VSS.n923 150
R4122 VSS.n933 VSS.n932 150
R4123 VSS.n944 VSS.n943 150
R4124 VSS.n948 VSS.n947 150
R4125 VSS.n952 VSS.n951 150
R4126 VSS.n956 VSS.n955 150
R4127 VSS.n5137 VSS.n5136 150
R4128 VSS.n441 VSS.n440 150
R4129 VSS.n5124 VSS.n439 150
R4130 VSS.n864 VSS.n863 150
R4131 VSS.n529 VSS.n528 150
R4132 VSS.n525 VSS.n524 150
R4133 VSS.n521 VSS.n520 150
R4134 VSS.n517 VSS.n516 150
R4135 VSS.n5103 VSS.n489 150
R4136 VSS.n5071 VSS.n5070 150
R4137 VSS.n710 VSS.n709 150
R4138 VSS.n5058 VSS.n5057 150
R4139 VSS.n695 VSS.n694 150
R4140 VSS.n691 VSS.n690 150
R4141 VSS.n687 VSS.n686 150
R4142 VSS.n683 VSS.n682 150
R4143 VSS.n5118 VSS.n5117 150
R4144 VSS.n472 VSS.n471 150
R4145 VSS.n5105 VSS.n470 150
R4146 VSS.n914 VSS.n478 150
R4147 VSS.n910 VSS.n478 150
R4148 VSS.n896 VSS.n895 150
R4149 VSS.n900 VSS.n899 150
R4150 VSS.n904 VSS.n903 150
R4151 VSS.n908 VSS.n907 150
R4152 VSS.n4570 VSS.n4527 150
R4153 VSS.n4568 VSS.n4528 150
R4154 VSS.n4555 VSS.n4542 150
R4155 VSS.n4553 VSS.n30 150
R4156 VSS.n4522 VSS.n4508 150
R4157 VSS.n4518 VSS.n4516 150
R4158 VSS.n4514 VSS.n4511 150
R4159 VSS.n5481 VSS.n55 150
R4160 VSS.n5487 VSS.n5483 150
R4161 VSS.n5487 VSS.n5486 150
R4162 VSS.n5499 VSS.n46 150
R4163 VSS.n5502 VSS.n5501 150
R4164 VSS.n5504 VSS.n43 150
R4165 VSS.n5527 VSS.n5526 150
R4166 VSS.n5524 VSS.n32 150
R4167 VSS.n5520 VSS.n5519 150
R4168 VSS.n5517 VSS.n35 150
R4169 VSS.n1695 VSS.n1694 150
R4170 VSS.n4367 VSS.n4366 150
R4171 VSS.n1721 VSS.n1720 150
R4172 VSS.n1726 VSS.n1411 150
R4173 VSS.n4581 VSS.n1410 150
R4174 VSS.n1424 VSS.n1423 150
R4175 VSS.n1428 VSS.n1427 150
R4176 VSS.n1432 VSS.n1421 150
R4177 VSS.n4578 VSS.n1443 150
R4178 VSS.n4565 VSS.n4564 150
R4179 VSS.n4537 VSS.n4536 150
R4180 VSS.n4550 VSS.n4549 150
R4181 VSS.n4392 VSS.n4391 150
R4182 VSS.n4388 VSS.n4387 150
R4183 VSS.n4384 VSS.n4383 150
R4184 VSS.n4380 VSS.n1442 150
R4185 VSS.n1756 VSS.n1749 150
R4186 VSS.n4346 VSS.n4345 150
R4187 VSS.n2425 VSS.n2424 150
R4188 VSS.n2433 VSS.n2432 150
R4189 VSS.n2407 VSS.n2406 150
R4190 VSS.n2403 VSS.n2402 150
R4191 VSS.n2399 VSS.n2398 150
R4192 VSS.n2395 VSS.n2394 150
R4193 VSS.n4378 VSS.n4377 150
R4194 VSS.n1705 VSS.n1704 150
R4195 VSS.n4363 VSS.n1702 150
R4196 VSS.n1724 VSS.n1723 150
R4197 VSS.n4312 VSS.n4311 150
R4198 VSS.n4308 VSS.n4307 150
R4199 VSS.n4304 VSS.n4303 150
R4200 VSS.n4300 VSS.n4299 150
R4201 VSS.n3672 VSS.n3485 150
R4202 VSS.n3520 VSS.n3515 150
R4203 VSS.n3561 VSS.n3516 150
R4204 VSS.n3547 VSS.n3491 150
R4205 VSS.n3500 VSS.n3499 150
R4206 VSS.n3504 VSS.n3503 150
R4207 VSS.n3508 VSS.n3507 150
R4208 VSS.n3512 VSS.n3497 150
R4209 VSS.n3669 VSS.n3488 150
R4210 VSS.n3633 VSS.n3488 150
R4211 VSS.n3659 VSS.n3658 150
R4212 VSS.n3642 VSS.n3641 150
R4213 VSS.n3648 VSS.n3647 150
R4214 VSS.n3609 VSS.n3608 150
R4215 VSS.n3613 VSS.n3612 150
R4216 VSS.n3617 VSS.n3616 150
R4217 VSS.n3619 VSS.n3569 150
R4218 VSS.n1480 VSS.n1473 150
R4219 VSS.n4483 VSS.n4482 150
R4220 VSS.n1633 VSS.n1632 150
R4221 VSS.n1642 VSS.n1641 150
R4222 VSS.n1617 VSS.n1616 150
R4223 VSS.n1613 VSS.n1612 150
R4224 VSS.n1609 VSS.n1608 150
R4225 VSS.n1605 VSS.n1604 150
R4226 VSS.n3483 VSS.n3482 150
R4227 VSS.n3530 VSS.n3529 150
R4228 VSS.n3558 VSS.n3557 150
R4229 VSS.n3537 VSS.n1457 150
R4230 VSS.n3590 VSS.n3589 150
R4231 VSS.n3594 VSS.n3593 150
R4232 VSS.n3598 VSS.n3597 150
R4233 VSS.n3602 VSS.n3601 150
R4234 VSS.n4477 VSS.n1509 150
R4235 VSS.n4445 VSS.n4444 150
R4236 VSS.n1547 VSS.n1546 150
R4237 VSS.n4432 VSS.n4431 150
R4238 VSS.n3572 VSS.n3571 150
R4239 VSS.n3576 VSS.n3575 150
R4240 VSS.n3580 VSS.n3579 150
R4241 VSS.n3584 VSS.n3583 150
R4242 VSS.n4492 VSS.n4491 150
R4243 VSS.n1492 VSS.n1491 150
R4244 VSS.n4479 VSS.n1490 150
R4245 VSS.n1623 VSS.n1498 150
R4246 VSS.n1619 VSS.n1498 150
R4247 VSS.n1590 VSS.n1589 150
R4248 VSS.n1594 VSS.n1593 150
R4249 VSS.n1598 VSS.n1597 150
R4250 VSS.n1602 VSS.n1601 150
R4251 VSS.n844 VSS.n843 150
R4252 VSS.n4875 VSS.n4874 150
R4253 VSS.n3461 VSS.n3460 150
R4254 VSS.n3452 VSS.n822 150
R4255 VSS.n3445 VSS.n3444 150
R4256 VSS.n3441 VSS.n3440 150
R4257 VSS.n3437 VSS.n3436 150
R4258 VSS.n3433 VSS.n818 150
R4259 VSS.n4947 VSS.n819 150
R4260 VSS.n4916 VSS.n819 150
R4261 VSS.n4937 VSS.n4936 150
R4262 VSS.n4925 VSS.n4924 150
R4263 VSS.n4950 VSS.n817 150
R4264 VSS.n4892 VSS.n4891 150
R4265 VSS.n4896 VSS.n4895 150
R4266 VSS.n4900 VSS.n4899 150
R4267 VSS.n4902 VSS.n836 150
R4268 VSS.n1001 VSS.n994 150
R4269 VSS.n4856 VSS.n4855 150
R4270 VSS.n3719 VSS.n3718 150
R4271 VSS.n3728 VSS.n3727 150
R4272 VSS.n3703 VSS.n3702 150
R4273 VSS.n3699 VSS.n3698 150
R4274 VSS.n3695 VSS.n3694 150
R4275 VSS.n3691 VSS.n3690 150
R4276 VSS.n4884 VSS.n4883 150
R4277 VSS.n979 VSS.n978 150
R4278 VSS.n4871 VSS.n977 150
R4279 VSS.n3471 VSS.n3470 150
R4280 VSS.n4808 VSS.n4807 150
R4281 VSS.n4804 VSS.n4803 150
R4282 VSS.n4800 VSS.n4799 150
R4283 VSS.n4796 VSS.n4795 150
R4284 VSS.n4850 VSS.n1030 150
R4285 VSS.n3781 VSS.n3780 150
R4286 VSS.n3789 VSS.n3788 150
R4287 VSS.n3797 VSS.n3796 150
R4288 VSS.n4826 VSS.n4825 150
R4289 VSS.n4822 VSS.n4821 150
R4290 VSS.n4818 VSS.n4817 150
R4291 VSS.n4814 VSS.n4813 150
R4292 VSS.n4865 VSS.n4864 150
R4293 VSS.n1013 VSS.n1012 150
R4294 VSS.n4852 VSS.n1011 150
R4295 VSS.n3709 VSS.n1019 150
R4296 VSS.n3705 VSS.n1019 150
R4297 VSS.n3751 VSS.n3750 150
R4298 VSS.n3747 VSS.n3746 150
R4299 VSS.n3743 VSS.n3742 150
R4300 VSS.n3739 VSS.n3738 150
R4301 VSS.n2237 VSS.n2236 150
R4302 VSS.n2089 VSS.n2088 150
R4303 VSS.n2223 VSS.n2222 150
R4304 VSS.n2098 VSS.n249 150
R4305 VSS.n5304 VSS.n264 150
R4306 VSS.n5300 VSS.n5299 150
R4307 VSS.n5296 VSS.n5295 150
R4308 VSS.n5292 VSS.n5291 150
R4309 VSS.n5307 VSS.n5306 150
R4310 VSS.n5306 VSS.n244 150
R4311 VSS.n5274 VSS.n5273 150
R4312 VSS.n286 VSS.n285 150
R4313 VSS.n5261 VSS.n5260 150
R4314 VSS.n2202 VSS.n2201 150
R4315 VSS.n2198 VSS.n2197 150
R4316 VSS.n2194 VSS.n2193 150
R4317 VSS.n2190 VSS.n2189 150
R4318 VSS.n2738 VSS.n2737 150
R4319 VSS.n2740 VSS.n2071 150
R4320 VSS.n2144 VSS.n2142 150
R4321 VSS.n2166 VSS.n2123 150
R4322 VSS.n2734 VSS.n2073 150
R4323 VSS.n2730 VSS.n2728 150
R4324 VSS.n2726 VSS.n2075 150
R4325 VSS.n2722 VSS.n2720 150
R4326 VSS.n2718 VSS.n2077 150
R4327 VSS.n2233 VSS.n2231 150
R4328 VSS.n2217 VSS.n2216 150
R4329 VSS.n2219 VSS.n2214 150
R4330 VSS.n2214 VSS.n2097 150
R4331 VSS.n2174 VSS.n2103 150
R4332 VSS.n2178 VSS.n2176 150
R4333 VSS.n2182 VSS.n2101 150
R4334 VSS.n2186 VSS.n2184 150
R4335 VSS.n3015 VSS.n3014 150
R4336 VSS.n2866 VSS.n2865 150
R4337 VSS.n3001 VSS.n3000 150
R4338 VSS.n2875 VSS.n498 150
R4339 VSS.n5097 VSS.n513 150
R4340 VSS.n5093 VSS.n5092 150
R4341 VSS.n5089 VSS.n5088 150
R4342 VSS.n5085 VSS.n5084 150
R4343 VSS.n5100 VSS.n5099 150
R4344 VSS.n5099 VSS.n493 150
R4345 VSS.n5067 VSS.n5066 150
R4346 VSS.n714 VSS.n713 150
R4347 VSS.n5054 VSS.n5053 150
R4348 VSS.n2981 VSS.n2980 150
R4349 VSS.n2977 VSS.n2976 150
R4350 VSS.n2973 VSS.n2972 150
R4351 VSS.n2969 VSS.n2968 150
R4352 VSS.n3044 VSS.n3043 150
R4353 VSS.n3046 VSS.n2028 150
R4354 VSS.n2923 VSS.n2921 150
R4355 VSS.n2945 VSS.n2902 150
R4356 VSS.n3040 VSS.n2850 150
R4357 VSS.n3036 VSS.n3034 150
R4358 VSS.n3032 VSS.n2852 150
R4359 VSS.n3028 VSS.n3026 150
R4360 VSS.n3024 VSS.n2854 150
R4361 VSS.n3011 VSS.n3009 150
R4362 VSS.n2995 VSS.n2994 150
R4363 VSS.n2997 VSS.n2992 150
R4364 VSS.n2992 VSS.n2874 150
R4365 VSS.n2953 VSS.n2882 150
R4366 VSS.n2957 VSS.n2955 150
R4367 VSS.n2961 VSS.n2880 150
R4368 VSS.n2965 VSS.n2963 150
R4369 VSS.n3412 VSS.n3411 150
R4370 VSS.n3289 VSS.n3288 150
R4371 VSS.n3398 VSS.n3397 150
R4372 VSS.n3298 VSS.n1518 150
R4373 VSS.n4471 VSS.n1533 150
R4374 VSS.n4467 VSS.n4466 150
R4375 VSS.n4463 VSS.n4462 150
R4376 VSS.n4459 VSS.n4458 150
R4377 VSS.n4474 VSS.n4473 150
R4378 VSS.n4473 VSS.n1513 150
R4379 VSS.n4441 VSS.n4440 150
R4380 VSS.n1551 VSS.n1550 150
R4381 VSS.n4428 VSS.n4427 150
R4382 VSS.n3378 VSS.n3377 150
R4383 VSS.n3374 VSS.n3373 150
R4384 VSS.n3370 VSS.n3369 150
R4385 VSS.n3366 VSS.n3365 150
R4386 VSS.n3952 VSS.n3951 150
R4387 VSS.n3954 VSS.n1952 150
R4388 VSS.n3326 VSS.n3324 150
R4389 VSS.n3342 VSS.n3306 150
R4390 VSS.n3948 VSS.n3273 150
R4391 VSS.n3944 VSS.n3942 150
R4392 VSS.n3940 VSS.n3275 150
R4393 VSS.n3936 VSS.n3934 150
R4394 VSS.n3932 VSS.n3277 150
R4395 VSS.n3408 VSS.n3406 150
R4396 VSS.n3392 VSS.n3391 150
R4397 VSS.n3394 VSS.n3389 150
R4398 VSS.n3389 VSS.n3297 150
R4399 VSS.n3350 VSS.n3305 150
R4400 VSS.n3354 VSS.n3352 150
R4401 VSS.n3358 VSS.n3303 150
R4402 VSS.n3362 VSS.n3360 150
R4403 VSS.n2631 VSS.n2630 150
R4404 VSS.n2647 VSS.n2646 150
R4405 VSS.n2637 VSS.n2636 150
R4406 VSS.n2750 VSS.n2044 150
R4407 VSS.n2107 VSS.n2106 150
R4408 VSS.n2111 VSS.n2110 150
R4409 VSS.n2115 VSS.n2114 150
R4410 VSS.n2119 VSS.n2118 150
R4411 VSS.n2748 VSS.n2046 150
R4412 VSS.n2069 VSS.n2046 150
R4413 VSS.n2138 VSS.n2137 150
R4414 VSS.n2148 VSS.n2147 150
R4415 VSS.n2163 VSS.n2162 150
R4416 VSS.n2662 VSS.n2661 150
R4417 VSS.n2666 VSS.n2665 150
R4418 VSS.n2670 VSS.n2669 150
R4419 VSS.n2672 VSS.n2063 150
R4420 VSS.n4623 VSS.n1399 147.339
R4421 VSS.n1374 VSS.n1371 145.082
R4422 VSS.n1377 VSS.n1374 144.706
R4423 VSS.t29 VSS.t76 141.204
R4424 VSS.t7 VSS.t13 136.665
R4425 VSS.n4617 VSS.n4616 132.815
R4426 VSS.n4629 VSS.n1399 131.463
R4427 VSS.n4668 VSS.t31 130.673
R4428 VSS.n2533 VSS.t40 130.673
R4429 VSS.n4610 VSS.t44 130.673
R4430 VSS.t42 VSS.n5548 130.673
R4431 VSS.n358 VSS.t44 129.871
R4432 VSS.n5251 VSS.t40 129.871
R4433 VSS.n5044 VSS.t40 129.871
R4434 VSS.n5007 VSS.t40 129.871
R4435 VSS.n4418 VSS.t40 129.871
R4436 VSS.n1227 VSS.t31 129.871
R4437 VSS.n1307 VSS.t31 129.871
R4438 VSS.n3871 VSS.t31 129.871
R4439 VSS.n4047 VSS.t31 129.871
R4440 VSS.t33 VSS.n4719 129.871
R4441 VSS.n4075 VSS.t38 129.871
R4442 VSS.n3096 VSS.t38 129.871
R4443 VSS.n3181 VSS.t38 129.871
R4444 VSS.n5224 VSS.t44 129
R4445 VSS.n5241 VSS.t40 129
R4446 VSS.n5034 VSS.t40 129
R4447 VSS.n4997 VSS.t40 129
R4448 VSS.n4408 VSS.t40 129
R4449 VSS.n1228 VSS.t31 129
R4450 VSS.n1306 VSS.t31 129
R4451 VSS.n3870 VSS.t31 129
R4452 VSS.n4039 VSS.t31 129
R4453 VSS.t33 VSS.n1186 129
R4454 VSS.n3992 VSS.t38 129
R4455 VSS.n3088 VSS.t38 129
R4456 VSS.n3177 VSS.t38 129
R4457 VSS.n4628 VSS.n4627 125.365
R4458 VSS.n4597 VSS.n21 124.832
R4459 VSS.n4643 VSS.n1386 124.832
R4460 VSS.n4192 VSS.n1359 124.832
R4461 VSS.n2707 VSS.n2571 124.832
R4462 VSS.t14 VSS.t28 120.034
R4463 VSS.n4634 VSS.n1395 117.469
R4464 VSS.n4638 VSS.n1394 116.469
R4465 VSS.n1358 VSS.n1185 115.677
R4466 VSS.t24 VSS.t63 115.597
R4467 VSS.t20 VSS.t24 115.597
R4468 VSS.t22 VSS.t20 115.597
R4469 VSS.t76 VSS.t22 115.597
R4470 VSS.n5564 VSS.n3 113.062
R4471 VSS.n4638 VSS.n4637 112.596
R4472 VSS.n1890 VSS.t29 110.477
R4473 VSS.n5565 VSS.n2 109.576
R4474 VSS.t11 VSS.t81 109.188
R4475 VSS.t3 VSS.t87 109.188
R4476 VSS.n1872 VSS.t16 107.017
R4477 VSS.n1397 VSS.n1395 106.951
R4478 VSS.n1889 VSS.t78 105.88
R4479 VSS.n2789 VSS.n2034 103.938
R4480 VSS.n1896 VSS.n1895 100.096
R4481 VSS.n1881 VSS.n1880 100.088
R4482 VSS.n1891 VSS.t35 99.5017
R4483 VSS.n5235 VSS.n322 98.5005
R4484 VSS.n5233 VSS.n329 98.5005
R4485 VSS.n760 VSS.n328 98.5005
R4486 VSS.n1584 VSS.n327 98.5005
R4487 VSS.n4643 VSS.n1389 98.5005
R4488 VSS.n5435 VSS.n80 98.5005
R4489 VSS.n965 VSS.n79 98.5005
R4490 VSS.n3681 VSS.n78 98.5005
R4491 VSS.n3540 VSS.n72 98.5005
R4492 VSS.n5535 VSS.n21 98.5005
R4493 VSS.n5255 VSS.n296 98.5005
R4494 VSS.n5048 VSS.n724 98.5005
R4495 VSS.n5010 VSS.n735 98.5005
R4496 VSS.n4422 VSS.n734 98.5005
R4497 VSS.n2514 VSS.n2392 98.5005
R4498 VSS.n4685 VSS.n1221 98.5005
R4499 VSS.n1341 VSS.n1276 98.5005
R4500 VSS.n3922 VSS.n3921 98.5005
R4501 VSS.n4050 VSS.n4011 98.5005
R4502 VSS.n4681 VSS.n1359 98.5005
R4503 VSS.n4712 VSS.n1201 98.5005
R4504 VSS.n4714 VSS.n1197 98.5005
R4505 VSS.n4734 VSS.n1158 98.5005
R4506 VSS.n3970 VSS.n1200 98.5005
R4507 VSS.n4214 VSS.n1850 98.5005
R4508 VSS.n2757 VSS.n2035 97.5252
R4509 VSS.n5422 VSS.n98 97.5252
R4510 VSS.n5209 VSS.n397 97.5252
R4511 VSS.n5470 VSS.n58 97.5252
R4512 VSS.n4956 VSS.n812 97.5252
R4513 VSS.n3063 VSS.n1992 97.5252
R4514 VSS.n3149 VSS.n1958 97.5252
R4515 VSS.n4077 VSS.n1912 97.5252
R4516 VSS.n2364 VSS.n2363 93.6243
R4517 VSS.n643 VSS.n320 93.6243
R4518 VSS.n5230 VSS.n324 93.6243
R4519 VSS.n4990 VSS.n325 93.6243
R4520 VSS.n4401 VSS.n326 93.6243
R4521 VSS.n2301 VSS.n2284 93.6243
R4522 VSS.n5432 VSS.n75 93.6243
R4523 VSS.n967 VSS.n76 93.6243
R4524 VSS.n3679 VSS.n77 93.6243
R4525 VSS.n5437 VSS.n73 93.6243
R4526 VSS.n5287 VSS.n268 93.6243
R4527 VSS.n5080 VSS.n698 93.6243
R4528 VSS.n5012 VSS.n731 93.6243
R4529 VSS.n4454 VSS.n732 93.6243
R4530 VSS.n4319 VSS.n733 93.6243
R4531 VSS.n2708 VSS.n2707 93.6243
R4532 VSS.n4688 VSS.n4687 93.6243
R4533 VSS.n1304 VSS.n1277 93.6243
R4534 VSS.n3919 VSS.n3868 93.6243
R4535 VSS.n4013 VSS.n4009 93.6243
R4536 VSS.n2681 VSS.n2677 93.6243
R4537 VSS.n2844 VSS.n1198 93.6243
R4538 VSS.n4766 VSS.n1130 93.6243
R4539 VSS.n3267 VSS.n1165 93.6243
R4540 VSS.n1836 VSS.n1199 93.6243
R4541 VSS.n5476 VSS.n58 89.7233
R4542 VSS.n5163 VSS.n98 89.7233
R4543 VSS.n3627 VSS.n812 89.7233
R4544 VSS.n4910 VSS.n397 89.7233
R4545 VSS.n2793 VSS.n2035 89.7233
R4546 VSS.n3113 VSS.n1992 89.7233
R4547 VSS.n4079 VSS.n4077 89.7233
R4548 VSS.n3185 VSS.n1958 89.7233
R4549 VSS.n673 VSS.n645 87.7728
R4550 VSS.n673 VSS.n647 87.7728
R4551 VSS.n669 VSS.n647 87.7728
R4552 VSS.n669 VSS.n666 87.7728
R4553 VSS.n666 VSS.n665 87.7728
R4554 VSS.n665 VSS.n649 87.7728
R4555 VSS.n661 VSS.n649 87.7728
R4556 VSS.n661 VSS.n652 87.7728
R4557 VSS.n657 VSS.n652 87.7728
R4558 VSS.n657 VSS.n654 87.7728
R4559 VSS.n5223 VSS.n342 87.7728
R4560 VSS.n4984 VSS.n765 87.7728
R4561 VSS.n4984 VSS.n767 87.7728
R4562 VSS.n4980 VSS.n767 87.7728
R4563 VSS.n4980 VSS.n4977 87.7728
R4564 VSS.n4977 VSS.n4976 87.7728
R4565 VSS.n4976 VSS.n769 87.7728
R4566 VSS.n4972 VSS.n769 87.7728
R4567 VSS.n4972 VSS.n772 87.7728
R4568 VSS.n4968 VSS.n772 87.7728
R4569 VSS.n4968 VSS.n4965 87.7728
R4570 VSS.n1682 VSS.n1654 87.7728
R4571 VSS.n1682 VSS.n1656 87.7728
R4572 VSS.n1678 VSS.n1656 87.7728
R4573 VSS.n1678 VSS.n1675 87.7728
R4574 VSS.n1675 VSS.n1674 87.7728
R4575 VSS.n1674 VSS.n1658 87.7728
R4576 VSS.n1670 VSS.n1658 87.7728
R4577 VSS.n1670 VSS.n1661 87.7728
R4578 VSS.n1666 VSS.n1661 87.7728
R4579 VSS.n1666 VSS.n71 87.7728
R4580 VSS.n4705 VSS.n1208 87.7728
R4581 VSS.n4705 VSS.n4704 87.7728
R4582 VSS.n4704 VSS.n1212 87.7728
R4583 VSS.n4700 VSS.n1212 87.7728
R4584 VSS.n4700 VSS.n4699 87.7728
R4585 VSS.n4699 VSS.n4698 87.7728
R4586 VSS.n4698 VSS.n1214 87.7728
R4587 VSS.n4694 VSS.n1214 87.7728
R4588 VSS.n4694 VSS.n1217 87.7728
R4589 VSS.n4690 VSS.n1217 87.7728
R4590 VSS.n4726 VSS.n1163 87.7728
R4591 VSS.n4726 VSS.n4725 87.7728
R4592 VSS.n4725 VSS.n1168 87.7728
R4593 VSS.n4721 VSS.n1168 87.7728
R4594 VSS.n4721 VSS.n1170 87.7728
R4595 VSS.n3908 VSS.n1170 87.7728
R4596 VSS.n3912 VSS.n3908 87.7728
R4597 VSS.n3912 VSS.n3906 87.7728
R4598 VSS.n3916 VSS.n3906 87.7728
R4599 VSS.n3917 VSS.n3916 87.7728
R4600 VSS.n4069 VSS.n3999 87.7728
R4601 VSS.n4069 VSS.n4002 87.7728
R4602 VSS.n4065 VSS.n4002 87.7728
R4603 VSS.n4065 VSS.n4063 87.7728
R4604 VSS.n4063 VSS.n4062 87.7728
R4605 VSS.n4062 VSS.n4004 87.7728
R4606 VSS.n4058 VSS.n4004 87.7728
R4607 VSS.n4058 VSS.n4006 87.7728
R4608 VSS.n4054 VSS.n4006 87.7728
R4609 VSS.n4054 VSS.n4008 87.7728
R4610 VSS.n2786 VSS.n2037 87.7728
R4611 VSS.n2786 VSS.n2762 87.7728
R4612 VSS.n2782 VSS.n2762 87.7728
R4613 VSS.n2782 VSS.n2779 87.7728
R4614 VSS.n2779 VSS.n2778 87.7728
R4615 VSS.n2778 VSS.n2764 87.7728
R4616 VSS.n2774 VSS.n2764 87.7728
R4617 VSS.n2774 VSS.n2770 87.7728
R4618 VSS.n2770 VSS.n2769 87.7728
R4619 VSS.n2769 VSS.n1205 87.7728
R4620 VSS.t2 VSS.t89 87.4943
R4621 VSS.n1882 VSS.t64 87.478
R4622 VSS.t89 VSS.t12 81.7096
R4623 VSS.n3097 VSS.n1992 79.9708
R4624 VSS.n3182 VSS.n1958 79.9708
R4625 VSS.n4077 VSS.n4076 79.9708
R4626 VSS.n2790 VSS.n2035 79.9708
R4627 VSS.n1886 VSS.n1884 79.0663
R4628 VSS.n5566 VSS.n5565 78.9338
R4629 VSS.n1886 VSS.n1885 78.778
R4630 VSS.t79 VSS.t7 77.3711
R4631 VSS.n2542 VSS.n2541 76.3222
R4632 VSS.n1855 VSS.n1851 76.3222
R4633 VSS.n2267 VSS.n2265 76.3222
R4634 VSS.n2388 VSS.n2387 76.3222
R4635 VSS.n2676 VSS.n2582 76.3222
R4636 VSS.n2297 VSS.n2279 76.3222
R4637 VSS.n2621 VSS.n2590 76.3222
R4638 VSS.n4158 VSS.n4157 76.3222
R4639 VSS.n2621 VSS.n2620 76.3222
R4640 VSS.n2582 VSS.n2580 76.3222
R4641 VSS.n2387 VSS.n2386 76.3222
R4642 VSS.n2268 VSS.n2267 76.3222
R4643 VSS.n2297 VSS.n2296 76.3222
R4644 VSS.n4158 VSS.n1869 76.3222
R4645 VSS.n4181 VSS.n1851 76.3222
R4646 VSS.n2543 VSS.n2542 76.3222
R4647 VSS.n4271 VSS.n1803 76.062
R4648 VSS.n1808 VSS.n1803 76.062
R4649 VSS.n2479 VSS.n1767 74.5978
R4650 VSS.n933 VSS.n448 74.5978
R4651 VSS.n943 VSS.n448 74.5978
R4652 VSS.n4580 VSS.n1411 74.5978
R4653 VSS.n2433 VSS.n1741 74.5978
R4654 VSS.n4581 VSS.n4580 74.5978
R4655 VSS.n1642 VSS.n1464 74.5978
R4656 VSS.n1617 VSS.n1464 74.5978
R4657 VSS.n3728 VSS.n986 74.5978
R4658 VSS.n3703 VSS.n986 74.5978
R4659 VSS.n2492 VSS.n1767 74.5978
R4660 VSS.n2407 VSS.n1741 74.5978
R4661 VSS.n676 VSS.n675 72.8181
R4662 VSS.n4987 VSS.n4986 72.8181
R4663 VSS.n1685 VSS.n1684 72.8181
R4664 VSS.n4357 VSS.n1753 69.3109
R4665 VSS.n4276 VSS.n1812 69.3109
R4666 VSS.n4276 VSS.n4275 69.3109
R4667 VSS.n3963 VSS.n3962 69.3109
R4668 VSS.n3963 VSS.n1944 69.3109
R4669 VSS.n4776 VSS.n1090 69.3109
R4670 VSS.n4769 VSS.n1090 69.3109
R4671 VSS.n3055 VSS.n3054 69.3109
R4672 VSS.n3055 VSS.n2020 69.3109
R4673 VSS.n4847 VSS.n1033 69.3109
R4674 VSS.n4831 VSS.n1033 69.3109
R4675 VSS.n1081 VSS.n1080 69.3109
R4676 VSS.n1113 VSS.n1081 69.3109
R4677 VSS.n5327 VSS.n204 69.3109
R4678 VSS.n2354 VSS.n204 69.3109
R4679 VSS.n5414 VSS.n5413 69.3109
R4680 VSS.n5414 VSS.n122 69.3109
R4681 VSS.n5347 VSS.n171 69.3109
R4682 VSS.n2324 VSS.n171 69.3109
R4683 VSS.n5201 VSS.n5200 69.3109
R4684 VSS.n5137 VSS.n425 69.3109
R4685 VSS.n516 VSS.n425 69.3109
R4686 VSS.n5201 VSS.n421 69.3109
R4687 VSS.n5118 VSS.n460 69.3109
R4688 VSS.n682 VSS.n460 69.3109
R4689 VSS.n5483 VSS.n5482 69.3109
R4690 VSS.n5482 VSS.n5481 69.3109
R4691 VSS.n4579 VSS.n4578 69.3109
R4692 VSS.n4378 VSS.n1691 69.3109
R4693 VSS.n4299 VSS.n1691 69.3109
R4694 VSS.n4579 VSS.n1442 69.3109
R4695 VSS.n3670 VSS.n3669 69.3109
R4696 VSS.n3482 VSS.n1468 69.3109
R4697 VSS.n3602 VSS.n1468 69.3109
R4698 VSS.n3670 VSS.n3569 69.3109
R4699 VSS.n4492 VSS.n1477 69.3109
R4700 VSS.n3584 VSS.n1477 69.3109
R4701 VSS.n4948 VSS.n4947 69.3109
R4702 VSS.n4884 VSS.n840 69.3109
R4703 VSS.n4795 VSS.n840 69.3109
R4704 VSS.n4948 VSS.n836 69.3109
R4705 VSS.n4865 VSS.n998 69.3109
R4706 VSS.n4813 VSS.n998 69.3109
R4707 VSS.n5307 VSS.n243 69.3109
R4708 VSS.n5291 VSS.n243 69.3109
R4709 VSS.n2719 VSS.n2718 69.3109
R4710 VSS.n2720 VSS.n2719 69.3109
R4711 VSS.n5100 VSS.n492 69.3109
R4712 VSS.n5084 VSS.n492 69.3109
R4713 VSS.n3025 VSS.n3024 69.3109
R4714 VSS.n3026 VSS.n3025 69.3109
R4715 VSS.n4474 VSS.n1512 69.3109
R4716 VSS.n4458 VSS.n1512 69.3109
R4717 VSS.n3933 VSS.n3932 69.3109
R4718 VSS.n3934 VSS.n3933 69.3109
R4719 VSS.n2749 VSS.n2748 69.3109
R4720 VSS.n2749 VSS.n2063 69.3109
R4721 VSS.n4323 VSS.n1753 69.3109
R4722 VSS.n1893 VSS.t34 66.259
R4723 VSS.n1879 VSS.t66 66.2527
R4724 VSS.t51 VSS.n1795 65.8183
R4725 VSS.t51 VSS.n1796 65.8183
R4726 VSS.t51 VSS.n1797 65.8183
R4727 VSS.t51 VSS.n1798 65.8183
R4728 VSS.t60 VSS.n1817 65.8183
R4729 VSS.t60 VSS.n1818 65.8183
R4730 VSS.t60 VSS.n1819 65.8183
R4731 VSS.t60 VSS.n1820 65.8183
R4732 VSS.t60 VSS.n1827 65.8183
R4733 VSS.t60 VSS.n1828 65.8183
R4734 VSS.t60 VSS.n1829 65.8183
R4735 VSS.t60 VSS.n1830 65.8183
R4736 VSS.t47 VSS.n1931 65.8183
R4737 VSS.t47 VSS.n1932 65.8183
R4738 VSS.t47 VSS.n1933 65.8183
R4739 VSS.t47 VSS.n1934 65.8183
R4740 VSS.t47 VSS.n1940 65.8183
R4741 VSS.t47 VSS.n1941 65.8183
R4742 VSS.t47 VSS.n1942 65.8183
R4743 VSS.t47 VSS.n1943 65.8183
R4744 VSS.t71 VSS.n1097 65.8183
R4745 VSS.t71 VSS.n1098 65.8183
R4746 VSS.t71 VSS.n1099 65.8183
R4747 VSS.t71 VSS.n1100 65.8183
R4748 VSS.t71 VSS.n1107 65.8183
R4749 VSS.t71 VSS.n1108 65.8183
R4750 VSS.t71 VSS.n1109 65.8183
R4751 VSS.t71 VSS.n4774 65.8183
R4752 VSS.t74 VSS.n2006 65.8183
R4753 VSS.t74 VSS.n2007 65.8183
R4754 VSS.t74 VSS.n2008 65.8183
R4755 VSS.t74 VSS.n2009 65.8183
R4756 VSS.t74 VSS.n2016 65.8183
R4757 VSS.t74 VSS.n2017 65.8183
R4758 VSS.t74 VSS.n2018 65.8183
R4759 VSS.t74 VSS.n2019 65.8183
R4760 VSS.t61 VSS.n4845 65.8183
R4761 VSS.t61 VSS.n1052 65.8183
R4762 VSS.t61 VSS.n1051 65.8183
R4763 VSS.t61 VSS.n1050 65.8183
R4764 VSS.t50 VSS.n1082 65.8183
R4765 VSS.t50 VSS.n1083 65.8183
R4766 VSS.t50 VSS.n1084 65.8183
R4767 VSS.t50 VSS.n1085 65.8183
R4768 VSS.t50 VSS.n1079 65.8183
R4769 VSS.t50 VSS.n1078 65.8183
R4770 VSS.t50 VSS.n1077 65.8183
R4771 VSS.t50 VSS.n1076 65.8183
R4772 VSS.t61 VSS.n1040 65.8183
R4773 VSS.t61 VSS.n1041 65.8183
R4774 VSS.t61 VSS.n1042 65.8183
R4775 VSS.t61 VSS.n1043 65.8183
R4776 VSS.t39 VSS.n235 65.8183
R4777 VSS.t39 VSS.n236 65.8183
R4778 VSS.t39 VSS.n237 65.8183
R4779 VSS.t39 VSS.n238 65.8183
R4780 VSS.t39 VSS.n234 65.8183
R4781 VSS.t39 VSS.n233 65.8183
R4782 VSS.t39 VSS.n232 65.8183
R4783 VSS.t39 VSS.n231 65.8183
R4784 VSS.t41 VSS.n121 65.8183
R4785 VSS.t41 VSS.n120 65.8183
R4786 VSS.t41 VSS.n119 65.8183
R4787 VSS.t41 VSS.n118 65.8183
R4788 VSS.t72 VSS.n196 65.8183
R4789 VSS.t72 VSS.n197 65.8183
R4790 VSS.t72 VSS.n198 65.8183
R4791 VSS.t72 VSS.n199 65.8183
R4792 VSS.t72 VSS.n195 65.8183
R4793 VSS.t72 VSS.n194 65.8183
R4794 VSS.t72 VSS.n193 65.8183
R4795 VSS.t72 VSS.n192 65.8183
R4796 VSS.t41 VSS.n109 65.8183
R4797 VSS.t41 VSS.n110 65.8183
R4798 VSS.t41 VSS.n111 65.8183
R4799 VSS.t41 VSS.n112 65.8183
R4800 VSS.t41 VSS.n107 65.8183
R4801 VSS.t41 VSS.n114 65.8183
R4802 VSS.t41 VSS.n106 65.8183
R4803 VSS.t41 VSS.n117 65.8183
R4804 VSS.t72 VSS.n188 65.8183
R4805 VSS.n5331 VSS.t72 65.8183
R4806 VSS.t72 VSS.n172 65.8183
R4807 VSS.t72 VSS.n189 65.8183
R4808 VSS.t72 VSS.n187 65.8183
R4809 VSS.t72 VSS.n186 65.8183
R4810 VSS.t72 VSS.n185 65.8183
R4811 VSS.n5311 VSS.t39 65.8183
R4812 VSS.t39 VSS.n226 65.8183
R4813 VSS.t39 VSS.n205 65.8183
R4814 VSS.t53 VSS.n408 65.8183
R4815 VSS.t53 VSS.n409 65.8183
R4816 VSS.t53 VSS.n410 65.8183
R4817 VSS.t53 VSS.n411 65.8183
R4818 VSS.t43 VSS.n452 65.8183
R4819 VSS.t43 VSS.n453 65.8183
R4820 VSS.t43 VSS.n454 65.8183
R4821 VSS.t43 VSS.n455 65.8183
R4822 VSS.t53 VSS.n417 65.8183
R4823 VSS.t53 VSS.n418 65.8183
R4824 VSS.t53 VSS.n419 65.8183
R4825 VSS.t53 VSS.n420 65.8183
R4826 VSS.t53 VSS.n406 65.8183
R4827 VSS.t53 VSS.n413 65.8183
R4828 VSS.t53 VSS.n405 65.8183
R4829 VSS.t53 VSS.n416 65.8183
R4830 VSS.t43 VSS.n443 65.8183
R4831 VSS.t43 VSS.n442 65.8183
R4832 VSS.n5123 VSS.t43 65.8183
R4833 VSS.t43 VSS.n426 65.8183
R4834 VSS.t73 VSS.n484 65.8183
R4835 VSS.t73 VSS.n485 65.8183
R4836 VSS.t73 VSS.n486 65.8183
R4837 VSS.t73 VSS.n487 65.8183
R4838 VSS.t73 VSS.n483 65.8183
R4839 VSS.t73 VSS.n482 65.8183
R4840 VSS.t73 VSS.n481 65.8183
R4841 VSS.t73 VSS.n480 65.8183
R4842 VSS.t43 VSS.n447 65.8183
R4843 VSS.t43 VSS.n446 65.8183
R4844 VSS.t43 VSS.n445 65.8183
R4845 VSS.t43 VSS.n444 65.8183
R4846 VSS.n4523 VSS.t56 65.8183
R4847 VSS.n4517 VSS.t56 65.8183
R4848 VSS.n4515 VSS.t56 65.8183
R4849 VSS.n4510 VSS.t56 65.8183
R4850 VSS.t70 VSS.n1745 65.8183
R4851 VSS.t70 VSS.n1746 65.8183
R4852 VSS.t70 VSS.n1747 65.8183
R4853 VSS.t70 VSS.n1748 65.8183
R4854 VSS.t48 VSS.n1441 65.8183
R4855 VSS.t48 VSS.n1440 65.8183
R4856 VSS.t48 VSS.n1439 65.8183
R4857 VSS.t48 VSS.n1438 65.8183
R4858 VSS.t48 VSS.n1416 65.8183
R4859 VSS.t48 VSS.n1436 65.8183
R4860 VSS.t48 VSS.n1413 65.8183
R4861 VSS.t48 VSS.n1437 65.8183
R4862 VSS.t70 VSS.n1707 65.8183
R4863 VSS.t70 VSS.n1706 65.8183
R4864 VSS.n4362 VSS.t70 65.8183
R4865 VSS.t70 VSS.n1692 65.8183
R4866 VSS.t48 VSS.n1435 65.8183
R4867 VSS.t48 VSS.n1420 65.8183
R4868 VSS.t48 VSS.n1419 65.8183
R4869 VSS.t48 VSS.n1418 65.8183
R4870 VSS.n5518 VSS.t56 65.8183
R4871 VSS.n34 VSS.t56 65.8183
R4872 VSS.n5525 VSS.t56 65.8183
R4873 VSS.n5528 VSS.t56 65.8183
R4874 VSS.n4554 VSS.t56 65.8183
R4875 VSS.n4541 VSS.t56 65.8183
R4876 VSS.n4569 VSS.t56 65.8183
R4877 VSS.n4526 VSS.t56 65.8183
R4878 VSS.t48 VSS.n1417 65.8183
R4879 VSS.t48 VSS.n1415 65.8183
R4880 VSS.t48 VSS.n1414 65.8183
R4881 VSS.t48 VSS.n1412 65.8183
R4882 VSS.t54 VSS.n3492 65.8183
R4883 VSS.t54 VSS.n3493 65.8183
R4884 VSS.t54 VSS.n3494 65.8183
R4885 VSS.t54 VSS.n3496 65.8183
R4886 VSS.t45 VSS.n1469 65.8183
R4887 VSS.t45 VSS.n1470 65.8183
R4888 VSS.t45 VSS.n1471 65.8183
R4889 VSS.t45 VSS.n1472 65.8183
R4890 VSS.t54 VSS.n3565 65.8183
R4891 VSS.t54 VSS.n3566 65.8183
R4892 VSS.t54 VSS.n3567 65.8183
R4893 VSS.t54 VSS.n3568 65.8183
R4894 VSS.t54 VSS.n3490 65.8183
R4895 VSS.t54 VSS.n3562 65.8183
R4896 VSS.t54 VSS.n3489 65.8183
R4897 VSS.n3671 VSS.t54 65.8183
R4898 VSS.n4497 VSS.t45 65.8183
R4899 VSS.t45 VSS.n1460 65.8183
R4900 VSS.t45 VSS.n1459 65.8183
R4901 VSS.t45 VSS.n1458 65.8183
R4902 VSS.t49 VSS.n1504 65.8183
R4903 VSS.t49 VSS.n1505 65.8183
R4904 VSS.t49 VSS.n1506 65.8183
R4905 VSS.t49 VSS.n1507 65.8183
R4906 VSS.t49 VSS.n1503 65.8183
R4907 VSS.t49 VSS.n1502 65.8183
R4908 VSS.t49 VSS.n1501 65.8183
R4909 VSS.t49 VSS.n1500 65.8183
R4910 VSS.t45 VSS.n1455 65.8183
R4911 VSS.t45 VSS.n1463 65.8183
R4912 VSS.t45 VSS.n1462 65.8183
R4913 VSS.t45 VSS.n1461 65.8183
R4914 VSS.t45 VSS.n1465 65.8183
R4915 VSS.t45 VSS.n1466 65.8183
R4916 VSS.t45 VSS.n1467 65.8183
R4917 VSS.t45 VSS.n4496 65.8183
R4918 VSS.t49 VSS.n1496 65.8183
R4919 VSS.n4478 VSS.t49 65.8183
R4920 VSS.t49 VSS.n1478 65.8183
R4921 VSS.t65 VSS.n823 65.8183
R4922 VSS.t65 VSS.n824 65.8183
R4923 VSS.t65 VSS.n825 65.8183
R4924 VSS.t65 VSS.n826 65.8183
R4925 VSS.t55 VSS.n990 65.8183
R4926 VSS.t55 VSS.n991 65.8183
R4927 VSS.t55 VSS.n992 65.8183
R4928 VSS.t55 VSS.n993 65.8183
R4929 VSS.t65 VSS.n832 65.8183
R4930 VSS.t65 VSS.n833 65.8183
R4931 VSS.t65 VSS.n834 65.8183
R4932 VSS.t65 VSS.n835 65.8183
R4933 VSS.t65 VSS.n821 65.8183
R4934 VSS.t65 VSS.n828 65.8183
R4935 VSS.t65 VSS.n820 65.8183
R4936 VSS.t65 VSS.n831 65.8183
R4937 VSS.t55 VSS.n981 65.8183
R4938 VSS.t55 VSS.n980 65.8183
R4939 VSS.n4870 VSS.t55 65.8183
R4940 VSS.t55 VSS.n841 65.8183
R4941 VSS.t69 VSS.n1025 65.8183
R4942 VSS.t69 VSS.n1026 65.8183
R4943 VSS.t69 VSS.n1027 65.8183
R4944 VSS.t69 VSS.n1028 65.8183
R4945 VSS.t69 VSS.n1024 65.8183
R4946 VSS.t69 VSS.n1023 65.8183
R4947 VSS.t69 VSS.n1022 65.8183
R4948 VSS.t69 VSS.n1021 65.8183
R4949 VSS.t55 VSS.n985 65.8183
R4950 VSS.t55 VSS.n984 65.8183
R4951 VSS.t55 VSS.n983 65.8183
R4952 VSS.t55 VSS.n982 65.8183
R4953 VSS.t55 VSS.n987 65.8183
R4954 VSS.t55 VSS.n988 65.8183
R4955 VSS.t55 VSS.n989 65.8183
R4956 VSS.t55 VSS.n4869 65.8183
R4957 VSS.t69 VSS.n1017 65.8183
R4958 VSS.n4851 VSS.t69 65.8183
R4959 VSS.t69 VSS.n999 65.8183
R4960 VSS.t43 VSS.n449 65.8183
R4961 VSS.t43 VSS.n450 65.8183
R4962 VSS.t43 VSS.n451 65.8183
R4963 VSS.t43 VSS.n5122 65.8183
R4964 VSS.t73 VSS.n476 65.8183
R4965 VSS.n5104 VSS.t73 65.8183
R4966 VSS.t73 VSS.n461 65.8183
R4967 VSS.t30 VSS.n5305 65.8183
R4968 VSS.t30 VSS.n262 65.8183
R4969 VSS.t30 VSS.n261 65.8183
R4970 VSS.t30 VSS.n260 65.8183
R4971 VSS.n2735 VSS.t57 65.8183
R4972 VSS.n2729 VSS.t57 65.8183
R4973 VSS.n2727 VSS.t57 65.8183
R4974 VSS.n2721 VSS.t57 65.8183
R4975 VSS.n2183 VSS.t57 65.8183
R4976 VSS.n2177 VSS.t57 65.8183
R4977 VSS.n2175 VSS.t57 65.8183
R4978 VSS.n2169 VSS.t57 65.8183
R4979 VSS.t30 VSS.n250 65.8183
R4980 VSS.t30 VSS.n251 65.8183
R4981 VSS.t30 VSS.n252 65.8183
R4982 VSS.t30 VSS.n253 65.8183
R4983 VSS.t59 VSS.n5098 65.8183
R4984 VSS.t59 VSS.n511 65.8183
R4985 VSS.t59 VSS.n510 65.8183
R4986 VSS.t59 VSS.n509 65.8183
R4987 VSS.n3041 VSS.t52 65.8183
R4988 VSS.n3035 VSS.t52 65.8183
R4989 VSS.n3033 VSS.t52 65.8183
R4990 VSS.n3027 VSS.t52 65.8183
R4991 VSS.n2962 VSS.t52 65.8183
R4992 VSS.n2956 VSS.t52 65.8183
R4993 VSS.n2954 VSS.t52 65.8183
R4994 VSS.n2948 VSS.t52 65.8183
R4995 VSS.t59 VSS.n499 65.8183
R4996 VSS.t59 VSS.n500 65.8183
R4997 VSS.t59 VSS.n501 65.8183
R4998 VSS.t59 VSS.n502 65.8183
R4999 VSS.t59 VSS.n497 65.8183
R5000 VSS.t59 VSS.n505 65.8183
R5001 VSS.t59 VSS.n496 65.8183
R5002 VSS.t59 VSS.n508 65.8183
R5003 VSS.n2996 VSS.t52 65.8183
R5004 VSS.n2863 VSS.t52 65.8183
R5005 VSS.n3010 VSS.t52 65.8183
R5006 VSS.t30 VSS.n248 65.8183
R5007 VSS.t30 VSS.n256 65.8183
R5008 VSS.t30 VSS.n247 65.8183
R5009 VSS.t30 VSS.n259 65.8183
R5010 VSS.n2218 VSS.t57 65.8183
R5011 VSS.n2086 VSS.t57 65.8183
R5012 VSS.n2232 VSS.t57 65.8183
R5013 VSS.t46 VSS.n4472 65.8183
R5014 VSS.t46 VSS.n1531 65.8183
R5015 VSS.t46 VSS.n1530 65.8183
R5016 VSS.t46 VSS.n1529 65.8183
R5017 VSS.n3949 VSS.t32 65.8183
R5018 VSS.n3943 VSS.t32 65.8183
R5019 VSS.n3941 VSS.t32 65.8183
R5020 VSS.n3935 VSS.t32 65.8183
R5021 VSS.n3359 VSS.t32 65.8183
R5022 VSS.n3353 VSS.t32 65.8183
R5023 VSS.n3351 VSS.t32 65.8183
R5024 VSS.n3345 VSS.t32 65.8183
R5025 VSS.t46 VSS.n1519 65.8183
R5026 VSS.t46 VSS.n1520 65.8183
R5027 VSS.t46 VSS.n1521 65.8183
R5028 VSS.t46 VSS.n1522 65.8183
R5029 VSS.t46 VSS.n1517 65.8183
R5030 VSS.t46 VSS.n1525 65.8183
R5031 VSS.t46 VSS.n1516 65.8183
R5032 VSS.t46 VSS.n1528 65.8183
R5033 VSS.n3393 VSS.t32 65.8183
R5034 VSS.n3286 VSS.t32 65.8183
R5035 VSS.n3407 VSS.t32 65.8183
R5036 VSS.t61 VSS.n1038 65.8183
R5037 VSS.t61 VSS.n1046 65.8183
R5038 VSS.t61 VSS.n1037 65.8183
R5039 VSS.t61 VSS.n1049 65.8183
R5040 VSS.t50 VSS.n1072 65.8183
R5041 VSS.t50 VSS.n1070 65.8183
R5042 VSS.n4780 VSS.t50 65.8183
R5043 VSS.t37 VSS.n2049 65.8183
R5044 VSS.t37 VSS.n2050 65.8183
R5045 VSS.t37 VSS.n2051 65.8183
R5046 VSS.t37 VSS.n2052 65.8183
R5047 VSS.t37 VSS.n2059 65.8183
R5048 VSS.t37 VSS.n2060 65.8183
R5049 VSS.t37 VSS.n2061 65.8183
R5050 VSS.t37 VSS.n2062 65.8183
R5051 VSS.t37 VSS.n2048 65.8183
R5052 VSS.t37 VSS.n2055 65.8183
R5053 VSS.t37 VSS.n2047 65.8183
R5054 VSS.t37 VSS.n2058 65.8183
R5055 VSS.t74 VSS.n2005 65.8183
R5056 VSS.t74 VSS.n2012 65.8183
R5057 VSS.t74 VSS.n2004 65.8183
R5058 VSS.t74 VSS.n2015 65.8183
R5059 VSS.t71 VSS.n1095 65.8183
R5060 VSS.t71 VSS.n1103 65.8183
R5061 VSS.t71 VSS.n1094 65.8183
R5062 VSS.t71 VSS.n1106 65.8183
R5063 VSS.t47 VSS.n1929 65.8183
R5064 VSS.t47 VSS.n1936 65.8183
R5065 VSS.t47 VSS.n1928 65.8183
R5066 VSS.t47 VSS.n1939 65.8183
R5067 VSS.t60 VSS.n1815 65.8183
R5068 VSS.t60 VSS.n1823 65.8183
R5069 VSS.t60 VSS.n1814 65.8183
R5070 VSS.t60 VSS.n1826 65.8183
R5071 VSS.n2167 VSS.t57 65.8183
R5072 VSS.n2143 VSS.t57 65.8183
R5073 VSS.n2141 VSS.t57 65.8183
R5074 VSS.n2739 VSS.t57 65.8183
R5075 VSS.n2946 VSS.t52 65.8183
R5076 VSS.n2922 VSS.t52 65.8183
R5077 VSS.n2920 VSS.t52 65.8183
R5078 VSS.n3045 VSS.t52 65.8183
R5079 VSS.t50 VSS.n1073 65.8183
R5080 VSS.t50 VSS.n1071 65.8183
R5081 VSS.t50 VSS.n1069 65.8183
R5082 VSS.t50 VSS.n1068 65.8183
R5083 VSS.n3343 VSS.t32 65.8183
R5084 VSS.n3325 VSS.t32 65.8183
R5085 VSS.n3323 VSS.t32 65.8183
R5086 VSS.n3953 VSS.t32 65.8183
R5087 VSS.t51 VSS.n1793 65.8183
R5088 VSS.t51 VSS.n1801 65.8183
R5089 VSS.t51 VSS.n1792 65.8183
R5090 VSS.t37 VSS.n2054 65.8183
R5091 VSS.t37 VSS.n2056 65.8183
R5092 VSS.t37 VSS.n2057 65.8183
R5093 VSS.t74 VSS.n2011 65.8183
R5094 VSS.t74 VSS.n2013 65.8183
R5095 VSS.t74 VSS.n2014 65.8183
R5096 VSS.t71 VSS.n1102 65.8183
R5097 VSS.t71 VSS.n1104 65.8183
R5098 VSS.t71 VSS.n1105 65.8183
R5099 VSS.t47 VSS.n1935 65.8183
R5100 VSS.t47 VSS.n1937 65.8183
R5101 VSS.t47 VSS.n1938 65.8183
R5102 VSS.t60 VSS.n1822 65.8183
R5103 VSS.t60 VSS.n1824 65.8183
R5104 VSS.t60 VSS.n1825 65.8183
R5105 VSS.t51 VSS.n1804 65.8183
R5106 VSS.t51 VSS.n1805 65.8183
R5107 VSS.t51 VSS.n1806 65.8183
R5108 VSS.t51 VSS.n1807 65.8183
R5109 VSS.t58 VSS.n4337 65.8183
R5110 VSS.t58 VSS.n1776 65.8183
R5111 VSS.t58 VSS.n1775 65.8183
R5112 VSS.t58 VSS.n1774 65.8183
R5113 VSS.t58 VSS.n1765 65.8183
R5114 VSS.t58 VSS.n1772 65.8183
R5115 VSS.t58 VSS.n1763 65.8183
R5116 VSS.t58 VSS.n1773 65.8183
R5117 VSS.t51 VSS.n1800 65.8183
R5118 VSS.t51 VSS.n1802 65.8183
R5119 VSS.n4284 VSS.t51 65.8183
R5120 VSS.t51 VSS.n4283 65.8183
R5121 VSS.t58 VSS.n1771 65.8183
R5122 VSS.t58 VSS.n1770 65.8183
R5123 VSS.t58 VSS.n1769 65.8183
R5124 VSS.t58 VSS.n1768 65.8183
R5125 VSS.t70 VSS.n1740 65.8183
R5126 VSS.t70 VSS.n1710 65.8183
R5127 VSS.t70 VSS.n1709 65.8183
R5128 VSS.t70 VSS.n1708 65.8183
R5129 VSS.t39 VSS.n228 65.8183
R5130 VSS.t39 VSS.n227 65.8183
R5131 VSS.t39 VSS.n222 65.8183
R5132 VSS.t39 VSS.n221 65.8183
R5133 VSS.t73 VSS.n477 65.8183
R5134 VSS.t73 VSS.n475 65.8183
R5135 VSS.t73 VSS.n474 65.8183
R5136 VSS.t73 VSS.n473 65.8183
R5137 VSS.t69 VSS.n1018 65.8183
R5138 VSS.t69 VSS.n1016 65.8183
R5139 VSS.t69 VSS.n1015 65.8183
R5140 VSS.t69 VSS.n1014 65.8183
R5141 VSS.t49 VSS.n1497 65.8183
R5142 VSS.t49 VSS.n1495 65.8183
R5143 VSS.t49 VSS.n1494 65.8183
R5144 VSS.t49 VSS.n1493 65.8183
R5145 VSS.t70 VSS.n1742 65.8183
R5146 VSS.t70 VSS.n1743 65.8183
R5147 VSS.t70 VSS.n1744 65.8183
R5148 VSS.t70 VSS.n4361 65.8183
R5149 VSS.t30 VSS.n255 65.8183
R5150 VSS.t30 VSS.n257 65.8183
R5151 VSS.t30 VSS.n258 65.8183
R5152 VSS.t59 VSS.n504 65.8183
R5153 VSS.t59 VSS.n506 65.8183
R5154 VSS.t59 VSS.n507 65.8183
R5155 VSS.t61 VSS.n1045 65.8183
R5156 VSS.t61 VSS.n1047 65.8183
R5157 VSS.t61 VSS.n1048 65.8183
R5158 VSS.t46 VSS.n1524 65.8183
R5159 VSS.t46 VSS.n1526 65.8183
R5160 VSS.t46 VSS.n1527 65.8183
R5161 VSS.t58 VSS.n1766 65.8183
R5162 VSS.t58 VSS.n1764 65.8183
R5163 VSS.n4341 VSS.t58 65.8183
R5164 VSS.t58 VSS.n1754 65.8183
R5165 VSS.t41 VSS.n113 65.8183
R5166 VSS.t41 VSS.n115 65.8183
R5167 VSS.t41 VSS.n116 65.8183
R5168 VSS.t53 VSS.n412 65.8183
R5169 VSS.t53 VSS.n414 65.8183
R5170 VSS.t53 VSS.n415 65.8183
R5171 VSS.t65 VSS.n827 65.8183
R5172 VSS.t65 VSS.n829 65.8183
R5173 VSS.t65 VSS.n830 65.8183
R5174 VSS.t54 VSS.n3514 65.8183
R5175 VSS.t54 VSS.n3563 65.8183
R5176 VSS.t54 VSS.n3564 65.8183
R5177 VSS.n5503 VSS.t56 65.8183
R5178 VSS.n5500 VSS.t56 65.8183
R5179 VSS.n5484 VSS.t56 65.8183
R5180 VSS.t72 VSS.n191 64.1729
R5181 VSS.t39 VSS.n230 64.1729
R5182 VSS.t49 VSS.n1499 64.1729
R5183 VSS.t69 VSS.n1020 64.1729
R5184 VSS.t73 VSS.n479 64.1729
R5185 VSS.n2964 VSS.t52 64.1729
R5186 VSS.n2185 VSS.t57 64.1729
R5187 VSS.n3361 VSS.t32 64.1729
R5188 VSS.t50 VSS.n1075 64.1729
R5189 VSS.t37 VSS.n2053 64.1729
R5190 VSS.t74 VSS.n2010 64.1729
R5191 VSS.t71 VSS.n1101 64.1729
R5192 VSS.n3964 VSS.t47 64.1729
R5193 VSS.t60 VSS.n1821 64.1729
R5194 VSS.t51 VSS.n1799 64.1729
R5195 VSS.t30 VSS.n254 64.1729
R5196 VSS.t59 VSS.n503 64.1729
R5197 VSS.t61 VSS.n1044 64.1729
R5198 VSS.t46 VSS.n1523 64.1729
R5199 VSS.n5415 VSS.t41 64.1729
R5200 VSS.n5202 VSS.t53 64.1729
R5201 VSS.n4949 VSS.t65 64.1729
R5202 VSS.t54 VSS.n3513 64.1729
R5203 VSS.n42 VSS.t56 64.1729
R5204 VSS.n5538 VSS.n21 62.4163
R5205 VSS.n4643 VSS.n1388 62.4163
R5206 VSS.n2543 VSS.n2392 62.4163
R5207 VSS.n4678 VSS.n1359 62.4163
R5208 VSS.n4181 VSS.n1850 62.4163
R5209 VSS.n2364 VSS.n2265 62.4163
R5210 VSS.n2388 VSS.n268 62.4163
R5211 VSS.n2707 VSS.n2570 62.4163
R5212 VSS.n2677 VSS.n2676 62.4163
R5213 VSS.n2301 VSS.n2279 62.4163
R5214 VSS.n1653 VSS.n1567 62.4163
R5215 VSS.n323 VSS.n303 62.4163
R5216 VSS.n654 VSS.n81 62.4163
R5217 VSS.n5218 VSS.n5217 62.4163
R5218 VSS.n764 VSS.n743 62.4163
R5219 VSS.n4965 VSS.n4964 62.4163
R5220 VSS.n5438 VSS.n71 62.4163
R5221 VSS.n300 VSS.n298 62.4163
R5222 VSS.n4690 VSS.n4689 62.4163
R5223 VSS.n1305 VSS.n1192 62.4163
R5224 VSS.n728 VSS.n726 62.4163
R5225 VSS.n5014 VSS.n330 62.4163
R5226 VSS.n1564 VSS.n1562 62.4163
R5227 VSS.n3917 VSS.n3904 62.4163
R5228 VSS.n739 VSS.n736 62.4163
R5229 VSS.n1195 VSS.n1193 62.4163
R5230 VSS.n1166 VSS.n1160 62.4163
R5231 VSS.n4074 VSS.n3973 62.4163
R5232 VSS.n4049 VSS.n4008 62.4163
R5233 VSS.n1205 VSS.n1202 62.4163
R5234 VSS.n4665 VSS.t31 62.1232
R5235 VSS.n4608 VSS.t44 62.1232
R5236 VSS.n5549 VSS.t42 62.1232
R5237 VSS.t0 VSS.t11 60.0169
R5238 VSS.t87 VSS.t0 60.0169
R5239 VSS.n4617 VSS.n1403 59.981
R5240 VSS.t72 VSS.n171 57.8461
R5241 VSS.t39 VSS.n204 57.8461
R5242 VSS.t43 VSS.n425 57.8461
R5243 VSS.t70 VSS.n1691 57.8461
R5244 VSS.t48 VSS.n4579 57.8461
R5245 VSS.t45 VSS.n1468 57.8461
R5246 VSS.t49 VSS.n1477 57.8461
R5247 VSS.t55 VSS.n840 57.8461
R5248 VSS.t69 VSS.n998 57.8461
R5249 VSS.t73 VSS.n460 57.8461
R5250 VSS.n3025 VSS.t52 57.8461
R5251 VSS.n2719 VSS.t57 57.8461
R5252 VSS.n3933 VSS.t32 57.8461
R5253 VSS.t50 VSS.n1081 57.8461
R5254 VSS.t37 VSS.n2749 57.8461
R5255 VSS.t74 VSS.n3055 57.8461
R5256 VSS.t71 VSS.n1090 57.8461
R5257 VSS.t47 VSS.n3963 57.8461
R5258 VSS.t60 VSS.n4276 57.8461
R5259 VSS.t30 VSS.n243 57.8461
R5260 VSS.t59 VSS.n492 57.8461
R5261 VSS.t61 VSS.n1033 57.8461
R5262 VSS.t46 VSS.n1512 57.8461
R5263 VSS.t58 VSS.n1753 57.8461
R5264 VSS.t41 VSS.n5414 57.8461
R5265 VSS.t53 VSS.n5201 57.8461
R5266 VSS.t65 VSS.n4948 57.8461
R5267 VSS.t54 VSS.n3670 57.8461
R5268 VSS.n5482 VSS.t56 57.8461
R5269 VSS.n2487 VSS.n1799 56.6572
R5270 VSS.n2451 VSS.n1799 56.6572
R5271 VSS.n4219 VSS.n1821 56.6572
R5272 VSS.n4131 VSS.n1821 56.6572
R5273 VSS.n3965 VSS.n3964 56.6572
R5274 VSS.n3964 VSS.n1926 56.6572
R5275 VSS.n4739 VSS.n1101 56.6572
R5276 VSS.n1962 VSS.n1101 56.6572
R5277 VSS.n2941 VSS.n2010 56.6572
R5278 VSS.n2898 VSS.n2010 56.6572
R5279 VSS.n3799 VSS.n1044 56.6572
R5280 VSS.n3830 VSS.n1075 56.6572
R5281 VSS.n3431 VSS.n1075 56.6572
R5282 VSS.n3813 VSS.n1044 56.6572
R5283 VSS.n613 VSS.n230 56.6572
R5284 VSS.n549 VSS.n230 56.6572
R5285 VSS.n5416 VSS.n5415 56.6572
R5286 VSS.n567 VSS.n191 56.6572
R5287 VSS.n597 VSS.n191 56.6572
R5288 VSS.n5415 VSS.n104 56.6572
R5289 VSS.n5203 VSS.n5202 56.6572
R5290 VSS.n5202 VSS.n403 56.6572
R5291 VSS.n910 VSS.n479 56.6572
R5292 VSS.n908 VSS.n479 56.6572
R5293 VSS.n43 VSS.n42 56.6572
R5294 VSS.n42 VSS.n35 56.6572
R5295 VSS.n3647 VSS.n3513 56.6572
R5296 VSS.n3513 VSS.n3512 56.6572
R5297 VSS.n1619 VSS.n1499 56.6572
R5298 VSS.n1602 VSS.n1499 56.6572
R5299 VSS.n4950 VSS.n4949 56.6572
R5300 VSS.n4949 VSS.n818 56.6572
R5301 VSS.n3705 VSS.n1020 56.6572
R5302 VSS.n3738 VSS.n1020 56.6572
R5303 VSS.n5260 VSS.n254 56.6572
R5304 VSS.n2185 VSS.n2097 56.6572
R5305 VSS.n2186 VSS.n2185 56.6572
R5306 VSS.n2189 VSS.n254 56.6572
R5307 VSS.n5053 VSS.n503 56.6572
R5308 VSS.n2964 VSS.n2874 56.6572
R5309 VSS.n2965 VSS.n2964 56.6572
R5310 VSS.n2968 VSS.n503 56.6572
R5311 VSS.n4427 VSS.n1523 56.6572
R5312 VSS.n3361 VSS.n3297 56.6572
R5313 VSS.n3362 VSS.n3361 56.6572
R5314 VSS.n3365 VSS.n1523 56.6572
R5315 VSS.n2162 VSS.n2053 56.6572
R5316 VSS.n2119 VSS.n2053 56.6572
R5317 VSS.n5561 VSS.n5560 56.3995
R5318 VSS.n2521 VSS.n2520 56.3995
R5319 VSS.n2300 VSS.n2278 56.3995
R5320 VSS.n2366 VSS.n2365 56.3995
R5321 VSS.n2253 VSS.n2252 56.3995
R5322 VSS.n5369 VSS.n167 56.3995
R5323 VSS.n2598 VSS.n2583 56.3995
R5324 VSS.n4177 VSS.n1852 56.3995
R5325 VSS.n2677 VSS.n2583 56.3995
R5326 VSS.n2252 VSS.n268 56.3995
R5327 VSS.n2365 VSS.n2364 56.3995
R5328 VSS.n2301 VSS.n2300 56.3995
R5329 VSS.n167 VSS.n166 56.3995
R5330 VSS.n1852 VSS.n1850 56.3995
R5331 VSS.n2520 VSS.n2392 56.3995
R5332 VSS.n5562 VSS.n5561 56.3995
R5333 VSS.n4660 VSS.n1373 55.7181
R5334 VSS.n1400 VSS.n1373 55.7181
R5335 VSS.n2545 VSS.t8 55.6967
R5336 VSS.n211 VSS.t44 55.4806
R5337 VSS.t42 VSS.n25 55.4806
R5338 VSS.t40 VSS.n270 55.4806
R5339 VSS.t33 VSS.n1132 55.4806
R5340 VSS.n1060 VSS.t31 55.4806
R5341 VSS.n4580 VSS.t48 55.2026
R5342 VSS.t45 VSS.n1464 55.2026
R5343 VSS.t55 VSS.n986 55.2026
R5344 VSS.t43 VSS.n448 55.2026
R5345 VSS.t58 VSS.n1767 55.2026
R5346 VSS.t70 VSS.n1741 55.2026
R5347 VSS.n4661 VSS.n1372 54.5887
R5348 VSS.n4621 VSS.n1372 54.5887
R5349 VSS.t51 VSS.n1803 54.4705
R5350 VSS.n1781 VSS.n1773 53.3664
R5351 VSS.n4288 VSS.n1763 53.3664
R5352 VSS.n2463 VSS.n1772 53.3664
R5353 VSS.n2472 VSS.n1765 53.3664
R5354 VSS.n2496 VSS.n1768 53.3664
R5355 VSS.n2500 VSS.n1769 53.3664
R5356 VSS.n2504 VSS.n1770 53.3664
R5357 VSS.n2508 VSS.n1771 53.3664
R5358 VSS.n4356 VSS.n1754 53.3664
R5359 VSS.n4341 VSS.n4340 53.3664
R5360 VSS.n1764 VSS.n1762 53.3664
R5361 VSS.n2429 VSS.n1766 53.3664
R5362 VSS.n4337 VSS.n4336 53.3664
R5363 VSS.n1778 VSS.n1776 53.3664
R5364 VSS.n4331 VSS.n1775 53.3664
R5365 VSS.n4327 VSS.n1774 53.3664
R5366 VSS.n1809 VSS.n1792 53.3664
R5367 VSS.n4244 VSS.n1801 53.3664
R5368 VSS.n4232 VSS.n1793 53.3664
R5369 VSS.n4270 VSS.n1804 53.3664
R5370 VSS.n4266 VSS.n1805 53.3664
R5371 VSS.n4262 VSS.n1806 53.3664
R5372 VSS.n4258 VSS.n1807 53.3664
R5373 VSS.n4283 VSS.n4282 53.3664
R5374 VSS.n4285 VSS.n4284 53.3664
R5375 VSS.n2459 VSS.n1802 53.3664
R5376 VSS.n2455 VSS.n1800 53.3664
R5377 VSS.n2438 VSS.n1798 53.3664
R5378 VSS.n2442 VSS.n1797 53.3664
R5379 VSS.n2446 VSS.n1796 53.3664
R5380 VSS.n2450 VSS.n1795 53.3664
R5381 VSS.n2447 VSS.n1795 53.3664
R5382 VSS.n2443 VSS.n1796 53.3664
R5383 VSS.n2439 VSS.n1797 53.3664
R5384 VSS.n2435 VSS.n1798 53.3664
R5385 VSS.n4096 VSS.n1826 53.3664
R5386 VSS.n4099 VSS.n1814 53.3664
R5387 VSS.n4112 VSS.n1823 53.3664
R5388 VSS.n4115 VSS.n1815 53.3664
R5389 VSS.n4144 VSS.n1820 53.3664
R5390 VSS.n4140 VSS.n1819 53.3664
R5391 VSS.n4136 VSS.n1818 53.3664
R5392 VSS.n4132 VSS.n1817 53.3664
R5393 VSS.n4135 VSS.n1817 53.3664
R5394 VSS.n4139 VSS.n1818 53.3664
R5395 VSS.n4143 VSS.n1819 53.3664
R5396 VSS.n4146 VSS.n1820 53.3664
R5397 VSS.n1825 VSS.n1813 53.3664
R5398 VSS.n4240 VSS.n1824 53.3664
R5399 VSS.n4228 VSS.n1822 53.3664
R5400 VSS.n4092 VSS.n1827 53.3664
R5401 VSS.n4091 VSS.n1828 53.3664
R5402 VSS.n4087 VSS.n1829 53.3664
R5403 VSS.n4083 VSS.n1830 53.3664
R5404 VSS.n4095 VSS.n1827 53.3664
R5405 VSS.n4088 VSS.n1828 53.3664
R5406 VSS.n4084 VSS.n1829 53.3664
R5407 VSS.n1831 VSS.n1830 53.3664
R5408 VSS.n3249 VSS.n1939 53.3664
R5409 VSS.n3192 VSS.n1928 53.3664
R5410 VSS.n3238 VSS.n1936 53.3664
R5411 VSS.n3201 VSS.n1929 53.3664
R5412 VSS.n3216 VSS.n1934 53.3664
R5413 VSS.n3212 VSS.n1933 53.3664
R5414 VSS.n3208 VSS.n1932 53.3664
R5415 VSS.n3204 VSS.n1931 53.3664
R5416 VSS.n3207 VSS.n1931 53.3664
R5417 VSS.n3211 VSS.n1932 53.3664
R5418 VSS.n3215 VSS.n1933 53.3664
R5419 VSS.n3218 VSS.n1934 53.3664
R5420 VSS.n1950 VSS.n1938 53.3664
R5421 VSS.n3320 VSS.n1937 53.3664
R5422 VSS.n3330 VSS.n1935 53.3664
R5423 VSS.n3253 VSS.n1940 53.3664
R5424 VSS.n3254 VSS.n1941 53.3664
R5425 VSS.n3258 VSS.n1942 53.3664
R5426 VSS.n3262 VSS.n1943 53.3664
R5427 VSS.n3250 VSS.n1940 53.3664
R5428 VSS.n3257 VSS.n1941 53.3664
R5429 VSS.n3261 VSS.n1942 53.3664
R5430 VSS.n3264 VSS.n1943 53.3664
R5431 VSS.n3107 VSS.n1106 53.3664
R5432 VSS.n3121 VSS.n1094 53.3664
R5433 VSS.n3124 VSS.n1103 53.3664
R5434 VSS.n3137 VSS.n1095 53.3664
R5435 VSS.n1975 VSS.n1100 53.3664
R5436 VSS.n1971 VSS.n1099 53.3664
R5437 VSS.n1967 VSS.n1098 53.3664
R5438 VSS.n1963 VSS.n1097 53.3664
R5439 VSS.n1966 VSS.n1097 53.3664
R5440 VSS.n1970 VSS.n1098 53.3664
R5441 VSS.n1974 VSS.n1099 53.3664
R5442 VSS.n1977 VSS.n1100 53.3664
R5443 VSS.n1105 VSS.n1091 53.3664
R5444 VSS.n4752 VSS.n1104 53.3664
R5445 VSS.n1148 VSS.n1102 53.3664
R5446 VSS.n3105 VSS.n1107 53.3664
R5447 VSS.n3104 VSS.n1108 53.3664
R5448 VSS.n3100 VSS.n1109 53.3664
R5449 VSS.n4774 VSS.n4773 53.3664
R5450 VSS.n3108 VSS.n1107 53.3664
R5451 VSS.n3101 VSS.n1108 53.3664
R5452 VSS.n1111 VSS.n1109 53.3664
R5453 VSS.n4774 VSS.n1110 53.3664
R5454 VSS.n2826 VSS.n2015 53.3664
R5455 VSS.n2800 VSS.n2004 53.3664
R5456 VSS.n2815 VSS.n2012 53.3664
R5457 VSS.n2806 VSS.n2005 53.3664
R5458 VSS.n2885 VSS.n2009 53.3664
R5459 VSS.n2889 VSS.n2008 53.3664
R5460 VSS.n2893 VSS.n2007 53.3664
R5461 VSS.n2897 VSS.n2006 53.3664
R5462 VSS.n2894 VSS.n2006 53.3664
R5463 VSS.n2890 VSS.n2007 53.3664
R5464 VSS.n2886 VSS.n2008 53.3664
R5465 VSS.n2009 VSS.n2002 53.3664
R5466 VSS.n2026 VSS.n2014 53.3664
R5467 VSS.n2917 VSS.n2013 53.3664
R5468 VSS.n2927 VSS.n2011 53.3664
R5469 VSS.n2830 VSS.n2016 53.3664
R5470 VSS.n2831 VSS.n2017 53.3664
R5471 VSS.n2835 VSS.n2018 53.3664
R5472 VSS.n2839 VSS.n2019 53.3664
R5473 VSS.n2827 VSS.n2016 53.3664
R5474 VSS.n2834 VSS.n2017 53.3664
R5475 VSS.n2838 VSS.n2018 53.3664
R5476 VSS.n2841 VSS.n2019 53.3664
R5477 VSS.n1057 VSS.n1049 53.3664
R5478 VSS.n4784 VSS.n1037 53.3664
R5479 VSS.n3841 VSS.n1046 53.3664
R5480 VSS.n3850 VSS.n1038 53.3664
R5481 VSS.n4845 VSS.n4844 53.3664
R5482 VSS.n1054 VSS.n1052 53.3664
R5483 VSS.n4839 VSS.n1051 53.3664
R5484 VSS.n4835 VSS.n1050 53.3664
R5485 VSS.n4845 VSS.n1053 53.3664
R5486 VSS.n4840 VSS.n1052 53.3664
R5487 VSS.n4836 VSS.n1051 53.3664
R5488 VSS.n4832 VSS.n1050 53.3664
R5489 VSS.n1048 VSS.n1034 53.3664
R5490 VSS.n3785 VSS.n1047 53.3664
R5491 VSS.n3793 VSS.n1045 53.3664
R5492 VSS.n3826 VSS.n1043 53.3664
R5493 VSS.n3822 VSS.n1042 53.3664
R5494 VSS.n3818 VSS.n1041 53.3664
R5495 VSS.n3814 VSS.n1040 53.3664
R5496 VSS.n1087 VSS.n1068 53.3664
R5497 VSS.n4756 VSS.n1069 53.3664
R5498 VSS.n1144 VSS.n1071 53.3664
R5499 VSS.n4743 VSS.n1073 53.3664
R5500 VSS.n1126 VSS.n1082 53.3664
R5501 VSS.n1125 VSS.n1083 53.3664
R5502 VSS.n1121 VSS.n1084 53.3664
R5503 VSS.n1117 VSS.n1085 53.3664
R5504 VSS.n1086 VSS.n1082 53.3664
R5505 VSS.n1122 VSS.n1083 53.3664
R5506 VSS.n1118 VSS.n1084 53.3664
R5507 VSS.n1114 VSS.n1085 53.3664
R5508 VSS.n4780 VSS.n1067 53.3664
R5509 VSS.n1070 VSS.n1066 53.3664
R5510 VSS.n3836 VSS.n1072 53.3664
R5511 VSS.n3418 VSS.n1076 53.3664
R5512 VSS.n3422 VSS.n1077 53.3664
R5513 VSS.n3426 VSS.n1078 53.3664
R5514 VSS.n3430 VSS.n1079 53.3664
R5515 VSS.n3427 VSS.n1079 53.3664
R5516 VSS.n3423 VSS.n1078 53.3664
R5517 VSS.n3419 VSS.n1077 53.3664
R5518 VSS.n3415 VSS.n1076 53.3664
R5519 VSS.n3817 VSS.n1040 53.3664
R5520 VSS.n3821 VSS.n1041 53.3664
R5521 VSS.n3825 VSS.n1042 53.3664
R5522 VSS.n3828 VSS.n1043 53.3664
R5523 VSS.n240 VSS.n221 53.3664
R5524 VSS.n5277 VSS.n222 53.3664
R5525 VSS.n282 VSS.n227 53.3664
R5526 VSS.n5264 VSS.n228 53.3664
R5527 VSS.n2341 VSS.n235 53.3664
R5528 VSS.n2342 VSS.n236 53.3664
R5529 VSS.n2346 VSS.n237 53.3664
R5530 VSS.n2350 VSS.n238 53.3664
R5531 VSS.n239 VSS.n235 53.3664
R5532 VSS.n2345 VSS.n236 53.3664
R5533 VSS.n2349 VSS.n237 53.3664
R5534 VSS.n2353 VSS.n238 53.3664
R5535 VSS.n5326 VSS.n205 53.3664
R5536 VSS.n226 VSS.n225 53.3664
R5537 VSS.n5312 VSS.n5311 53.3664
R5538 VSS.n536 VSS.n231 53.3664
R5539 VSS.n540 VSS.n232 53.3664
R5540 VSS.n544 VSS.n233 53.3664
R5541 VSS.n548 VSS.n234 53.3664
R5542 VSS.n545 VSS.n234 53.3664
R5543 VSS.n541 VSS.n233 53.3664
R5544 VSS.n537 VSS.n232 53.3664
R5545 VSS.n533 VSS.n231 53.3664
R5546 VSS.n5350 VSS.n117 53.3664
R5547 VSS.n175 VSS.n106 53.3664
R5548 VSS.n5336 VSS.n114 53.3664
R5549 VSS.n578 VSS.n107 53.3664
R5550 VSS.n5354 VSS.n121 53.3664
R5551 VSS.n5355 VSS.n120 53.3664
R5552 VSS.n5359 VSS.n119 53.3664
R5553 VSS.n5363 VSS.n118 53.3664
R5554 VSS.n5351 VSS.n121 53.3664
R5555 VSS.n5358 VSS.n120 53.3664
R5556 VSS.n5362 VSS.n119 53.3664
R5557 VSS.n5365 VSS.n118 53.3664
R5558 VSS.n131 VSS.n116 53.3664
R5559 VSS.n5402 VSS.n115 53.3664
R5560 VSS.n5391 VSS.n113 53.3664
R5561 VSS.n563 VSS.n112 53.3664
R5562 VSS.n559 VSS.n111 53.3664
R5563 VSS.n555 VSS.n110 53.3664
R5564 VSS.n551 VSS.n109 53.3664
R5565 VSS.n201 VSS.n185 53.3664
R5566 VSS.n214 VSS.n186 53.3664
R5567 VSS.n5315 VSS.n187 53.3664
R5568 VSS.n626 VSS.n189 53.3664
R5569 VSS.n2337 VSS.n196 53.3664
R5570 VSS.n2336 VSS.n197 53.3664
R5571 VSS.n2332 VSS.n198 53.3664
R5572 VSS.n2328 VSS.n199 53.3664
R5573 VSS.n200 VSS.n196 53.3664
R5574 VSS.n2333 VSS.n197 53.3664
R5575 VSS.n2329 VSS.n198 53.3664
R5576 VSS.n2325 VSS.n199 53.3664
R5577 VSS.n5346 VSS.n172 53.3664
R5578 VSS.n5331 VSS.n184 53.3664
R5579 VSS.n188 VSS.n181 53.3664
R5580 VSS.n610 VSS.n192 53.3664
R5581 VSS.n606 VSS.n193 53.3664
R5582 VSS.n602 VSS.n194 53.3664
R5583 VSS.n598 VSS.n195 53.3664
R5584 VSS.n601 VSS.n195 53.3664
R5585 VSS.n605 VSS.n194 53.3664
R5586 VSS.n609 VSS.n193 53.3664
R5587 VSS.n629 VSS.n192 53.3664
R5588 VSS.n554 VSS.n109 53.3664
R5589 VSS.n558 VSS.n110 53.3664
R5590 VSS.n562 VSS.n111 53.3664
R5591 VSS.n565 VSS.n112 53.3664
R5592 VSS.n585 VSS.n107 53.3664
R5593 VSS.n577 VSS.n114 53.3664
R5594 VSS.n5335 VSS.n106 53.3664
R5595 VSS.n174 VSS.n117 53.3664
R5596 VSS.n570 VSS.n188 53.3664
R5597 VSS.n5332 VSS.n5331 53.3664
R5598 VSS.n183 VSS.n172 53.3664
R5599 VSS.n630 VSS.n189 53.3664
R5600 VSS.n625 VSS.n187 53.3664
R5601 VSS.n5316 VSS.n186 53.3664
R5602 VSS.n213 VSS.n185 53.3664
R5603 VSS.n5311 VSS.n220 53.3664
R5604 VSS.n226 VSS.n219 53.3664
R5605 VSS.n224 VSS.n205 53.3664
R5606 VSS.n5140 VSS.n416 53.3664
R5607 VSS.n429 VSS.n405 53.3664
R5608 VSS.n5127 VSS.n413 53.3664
R5609 VSS.n861 VSS.n406 53.3664
R5610 VSS.n887 VSS.n411 53.3664
R5611 VSS.n883 VSS.n410 53.3664
R5612 VSS.n879 VSS.n409 53.3664
R5613 VSS.n875 VSS.n408 53.3664
R5614 VSS.n878 VSS.n408 53.3664
R5615 VSS.n882 VSS.n409 53.3664
R5616 VSS.n886 VSS.n410 53.3664
R5617 VSS.n889 VSS.n411 53.3664
R5618 VSS.n5169 VSS.n415 53.3664
R5619 VSS.n5189 VSS.n414 53.3664
R5620 VSS.n5178 VSS.n412 53.3664
R5621 VSS.n5144 VSS.n417 53.3664
R5622 VSS.n5145 VSS.n418 53.3664
R5623 VSS.n5149 VSS.n419 53.3664
R5624 VSS.n5153 VSS.n420 53.3664
R5625 VSS.n5122 VSS.n5121 53.3664
R5626 VSS.n463 VSS.n451 53.3664
R5627 VSS.n5108 VSS.n450 53.3664
R5628 VSS.n924 VSS.n449 53.3664
R5629 VSS.n947 VSS.n444 53.3664
R5630 VSS.n951 VSS.n445 53.3664
R5631 VSS.n955 VSS.n446 53.3664
R5632 VSS.n959 VSS.n447 53.3664
R5633 VSS.n5136 VSS.n426 53.3664
R5634 VSS.n5123 VSS.n441 53.3664
R5635 VSS.n442 VSS.n439 53.3664
R5636 VSS.n863 VSS.n443 53.3664
R5637 VSS.n529 VSS.n452 53.3664
R5638 VSS.n528 VSS.n453 53.3664
R5639 VSS.n524 VSS.n454 53.3664
R5640 VSS.n520 VSS.n455 53.3664
R5641 VSS.n457 VSS.n452 53.3664
R5642 VSS.n525 VSS.n453 53.3664
R5643 VSS.n521 VSS.n454 53.3664
R5644 VSS.n517 VSS.n455 53.3664
R5645 VSS.n5141 VSS.n417 53.3664
R5646 VSS.n5148 VSS.n418 53.3664
R5647 VSS.n5152 VSS.n419 53.3664
R5648 VSS.n5155 VSS.n420 53.3664
R5649 VSS.n866 VSS.n406 53.3664
R5650 VSS.n860 VSS.n413 53.3664
R5651 VSS.n5128 VSS.n405 53.3664
R5652 VSS.n428 VSS.n416 53.3664
R5653 VSS.n958 VSS.n443 53.3664
R5654 VSS.n864 VSS.n442 53.3664
R5655 VSS.n5124 VSS.n5123 53.3664
R5656 VSS.n440 VSS.n426 53.3664
R5657 VSS.n489 VSS.n473 53.3664
R5658 VSS.n5070 VSS.n474 53.3664
R5659 VSS.n710 VSS.n475 53.3664
R5660 VSS.n5057 VSS.n477 53.3664
R5661 VSS.n695 VSS.n484 53.3664
R5662 VSS.n694 VSS.n485 53.3664
R5663 VSS.n690 VSS.n486 53.3664
R5664 VSS.n686 VSS.n487 53.3664
R5665 VSS.n488 VSS.n484 53.3664
R5666 VSS.n691 VSS.n485 53.3664
R5667 VSS.n687 VSS.n486 53.3664
R5668 VSS.n683 VSS.n487 53.3664
R5669 VSS.n5117 VSS.n461 53.3664
R5670 VSS.n5104 VSS.n472 53.3664
R5671 VSS.n476 VSS.n470 53.3664
R5672 VSS.n895 VSS.n480 53.3664
R5673 VSS.n899 VSS.n481 53.3664
R5674 VSS.n903 VSS.n482 53.3664
R5675 VSS.n907 VSS.n483 53.3664
R5676 VSS.n904 VSS.n483 53.3664
R5677 VSS.n900 VSS.n482 53.3664
R5678 VSS.n896 VSS.n481 53.3664
R5679 VSS.n892 VSS.n480 53.3664
R5680 VSS.n956 VSS.n447 53.3664
R5681 VSS.n952 VSS.n446 53.3664
R5682 VSS.n948 VSS.n445 53.3664
R5683 VSS.n944 VSS.n444 53.3664
R5684 VSS.n4526 VSS.n4525 53.3664
R5685 VSS.n4570 VSS.n4569 53.3664
R5686 VSS.n4541 VSS.n4528 53.3664
R5687 VSS.n4555 VSS.n4554 53.3664
R5688 VSS.n4523 VSS.n4522 53.3664
R5689 VSS.n4517 VSS.n4508 53.3664
R5690 VSS.n4516 VSS.n4515 53.3664
R5691 VSS.n4511 VSS.n4510 53.3664
R5692 VSS.n4524 VSS.n4523 53.3664
R5693 VSS.n4518 VSS.n4517 53.3664
R5694 VSS.n4515 VSS.n4514 53.3664
R5695 VSS.n4510 VSS.n55 53.3664
R5696 VSS.n5486 VSS.n5484 53.3664
R5697 VSS.n5500 VSS.n5499 53.3664
R5698 VSS.n5503 VSS.n5502 53.3664
R5699 VSS.n5528 VSS.n5527 53.3664
R5700 VSS.n5525 VSS.n5524 53.3664
R5701 VSS.n5520 VSS.n34 53.3664
R5702 VSS.n5518 VSS.n5517 53.3664
R5703 VSS.n4396 VSS.n1437 53.3664
R5704 VSS.n1695 VSS.n1413 53.3664
R5705 VSS.n4367 VSS.n1436 53.3664
R5706 VSS.n1721 VSS.n1416 53.3664
R5707 VSS.n1423 VSS.n1418 53.3664
R5708 VSS.n1427 VSS.n1419 53.3664
R5709 VSS.n1421 VSS.n1420 53.3664
R5710 VSS.n1435 VSS.n1434 53.3664
R5711 VSS.n1443 VSS.n1412 53.3664
R5712 VSS.n4565 VSS.n1414 53.3664
R5713 VSS.n4537 VSS.n1415 53.3664
R5714 VSS.n4550 VSS.n1417 53.3664
R5715 VSS.n4392 VSS.n1441 53.3664
R5716 VSS.n4391 VSS.n1440 53.3664
R5717 VSS.n4387 VSS.n1439 53.3664
R5718 VSS.n4383 VSS.n1438 53.3664
R5719 VSS.n4361 VSS.n4360 53.3664
R5720 VSS.n1756 VSS.n1744 53.3664
R5721 VSS.n4346 VSS.n1743 53.3664
R5722 VSS.n2425 VSS.n1742 53.3664
R5723 VSS.n2403 VSS.n1708 53.3664
R5724 VSS.n2399 VSS.n1709 53.3664
R5725 VSS.n2395 VSS.n1710 53.3664
R5726 VSS.n1740 VSS.n1739 53.3664
R5727 VSS.n4377 VSS.n1692 53.3664
R5728 VSS.n4362 VSS.n1705 53.3664
R5729 VSS.n1706 VSS.n1702 53.3664
R5730 VSS.n1723 VSS.n1707 53.3664
R5731 VSS.n4312 VSS.n1745 53.3664
R5732 VSS.n4311 VSS.n1746 53.3664
R5733 VSS.n4307 VSS.n1747 53.3664
R5734 VSS.n4303 VSS.n1748 53.3664
R5735 VSS.n1750 VSS.n1745 53.3664
R5736 VSS.n4308 VSS.n1746 53.3664
R5737 VSS.n4304 VSS.n1747 53.3664
R5738 VSS.n4300 VSS.n1748 53.3664
R5739 VSS.n4395 VSS.n1441 53.3664
R5740 VSS.n4388 VSS.n1440 53.3664
R5741 VSS.n4384 VSS.n1439 53.3664
R5742 VSS.n4380 VSS.n1438 53.3664
R5743 VSS.n1726 VSS.n1416 53.3664
R5744 VSS.n1720 VSS.n1436 53.3664
R5745 VSS.n4366 VSS.n1413 53.3664
R5746 VSS.n1694 VSS.n1437 53.3664
R5747 VSS.n1738 VSS.n1707 53.3664
R5748 VSS.n1724 VSS.n1706 53.3664
R5749 VSS.n4363 VSS.n4362 53.3664
R5750 VSS.n1704 VSS.n1692 53.3664
R5751 VSS.n1435 VSS.n1432 53.3664
R5752 VSS.n1428 VSS.n1420 53.3664
R5753 VSS.n1424 VSS.n1419 53.3664
R5754 VSS.n1418 VSS.n1410 53.3664
R5755 VSS.n5519 VSS.n5518 53.3664
R5756 VSS.n34 VSS.n32 53.3664
R5757 VSS.n5526 VSS.n5525 53.3664
R5758 VSS.n5529 VSS.n5528 53.3664
R5759 VSS.n4554 VSS.n4553 53.3664
R5760 VSS.n4542 VSS.n4541 53.3664
R5761 VSS.n4569 VSS.n4568 53.3664
R5762 VSS.n4527 VSS.n4526 53.3664
R5763 VSS.n1433 VSS.n1417 53.3664
R5764 VSS.n4549 VSS.n1415 53.3664
R5765 VSS.n4536 VSS.n1414 53.3664
R5766 VSS.n4564 VSS.n1412 53.3664
R5767 VSS.n3671 VSS.n3487 53.3664
R5768 VSS.n3489 VSS.n3485 53.3664
R5769 VSS.n3562 VSS.n3515 53.3664
R5770 VSS.n3516 VSS.n3490 53.3664
R5771 VSS.n3499 VSS.n3496 53.3664
R5772 VSS.n3503 VSS.n3494 53.3664
R5773 VSS.n3507 VSS.n3493 53.3664
R5774 VSS.n3497 VSS.n3492 53.3664
R5775 VSS.n3508 VSS.n3492 53.3664
R5776 VSS.n3504 VSS.n3493 53.3664
R5777 VSS.n3500 VSS.n3494 53.3664
R5778 VSS.n3496 VSS.n3495 53.3664
R5779 VSS.n3633 VSS.n3564 53.3664
R5780 VSS.n3658 VSS.n3563 53.3664
R5781 VSS.n3642 VSS.n3514 53.3664
R5782 VSS.n3608 VSS.n3565 53.3664
R5783 VSS.n3609 VSS.n3566 53.3664
R5784 VSS.n3613 VSS.n3567 53.3664
R5785 VSS.n3617 VSS.n3568 53.3664
R5786 VSS.n4496 VSS.n4495 53.3664
R5787 VSS.n1480 VSS.n1467 53.3664
R5788 VSS.n4482 VSS.n1466 53.3664
R5789 VSS.n1633 VSS.n1465 53.3664
R5790 VSS.n1613 VSS.n1461 53.3664
R5791 VSS.n1609 VSS.n1462 53.3664
R5792 VSS.n1605 VSS.n1463 53.3664
R5793 VSS.n4499 VSS.n1455 53.3664
R5794 VSS.n3483 VSS.n1458 53.3664
R5795 VSS.n3530 VSS.n1459 53.3664
R5796 VSS.n3558 VSS.n1460 53.3664
R5797 VSS.n4497 VSS.n1457 53.3664
R5798 VSS.n3589 VSS.n1469 53.3664
R5799 VSS.n3590 VSS.n1470 53.3664
R5800 VSS.n3594 VSS.n1471 53.3664
R5801 VSS.n3598 VSS.n1472 53.3664
R5802 VSS.n1474 VSS.n1469 53.3664
R5803 VSS.n3593 VSS.n1470 53.3664
R5804 VSS.n3597 VSS.n1471 53.3664
R5805 VSS.n3601 VSS.n1472 53.3664
R5806 VSS.n3605 VSS.n3565 53.3664
R5807 VSS.n3612 VSS.n3566 53.3664
R5808 VSS.n3616 VSS.n3567 53.3664
R5809 VSS.n3619 VSS.n3568 53.3664
R5810 VSS.n3547 VSS.n3490 53.3664
R5811 VSS.n3562 VSS.n3561 53.3664
R5812 VSS.n3520 VSS.n3489 53.3664
R5813 VSS.n3672 VSS.n3671 53.3664
R5814 VSS.n4498 VSS.n4497 53.3664
R5815 VSS.n3537 VSS.n1460 53.3664
R5816 VSS.n3557 VSS.n1459 53.3664
R5817 VSS.n3529 VSS.n1458 53.3664
R5818 VSS.n1509 VSS.n1493 53.3664
R5819 VSS.n4444 VSS.n1494 53.3664
R5820 VSS.n1547 VSS.n1495 53.3664
R5821 VSS.n4431 VSS.n1497 53.3664
R5822 VSS.n3571 VSS.n1504 53.3664
R5823 VSS.n3572 VSS.n1505 53.3664
R5824 VSS.n3576 VSS.n1506 53.3664
R5825 VSS.n3580 VSS.n1507 53.3664
R5826 VSS.n1508 VSS.n1504 53.3664
R5827 VSS.n3575 VSS.n1505 53.3664
R5828 VSS.n3579 VSS.n1506 53.3664
R5829 VSS.n3583 VSS.n1507 53.3664
R5830 VSS.n4491 VSS.n1478 53.3664
R5831 VSS.n4478 VSS.n1492 53.3664
R5832 VSS.n1496 VSS.n1490 53.3664
R5833 VSS.n1589 VSS.n1500 53.3664
R5834 VSS.n1593 VSS.n1501 53.3664
R5835 VSS.n1597 VSS.n1502 53.3664
R5836 VSS.n1601 VSS.n1503 53.3664
R5837 VSS.n1598 VSS.n1503 53.3664
R5838 VSS.n1594 VSS.n1502 53.3664
R5839 VSS.n1590 VSS.n1501 53.3664
R5840 VSS.n1586 VSS.n1500 53.3664
R5841 VSS.n1604 VSS.n1455 53.3664
R5842 VSS.n1608 VSS.n1463 53.3664
R5843 VSS.n1612 VSS.n1462 53.3664
R5844 VSS.n1616 VSS.n1461 53.3664
R5845 VSS.n1641 VSS.n1465 53.3664
R5846 VSS.n1632 VSS.n1466 53.3664
R5847 VSS.n4483 VSS.n1467 53.3664
R5848 VSS.n4496 VSS.n1473 53.3664
R5849 VSS.n1623 VSS.n1496 53.3664
R5850 VSS.n4479 VSS.n4478 53.3664
R5851 VSS.n1491 VSS.n1478 53.3664
R5852 VSS.n4887 VSS.n831 53.3664
R5853 VSS.n844 VSS.n820 53.3664
R5854 VSS.n4874 VSS.n828 53.3664
R5855 VSS.n3460 VSS.n821 53.3664
R5856 VSS.n3445 VSS.n826 53.3664
R5857 VSS.n3441 VSS.n825 53.3664
R5858 VSS.n3437 VSS.n824 53.3664
R5859 VSS.n3433 VSS.n823 53.3664
R5860 VSS.n3436 VSS.n823 53.3664
R5861 VSS.n3440 VSS.n824 53.3664
R5862 VSS.n3444 VSS.n825 53.3664
R5863 VSS.n3447 VSS.n826 53.3664
R5864 VSS.n4916 VSS.n830 53.3664
R5865 VSS.n4936 VSS.n829 53.3664
R5866 VSS.n4925 VSS.n827 53.3664
R5867 VSS.n4891 VSS.n832 53.3664
R5868 VSS.n4892 VSS.n833 53.3664
R5869 VSS.n4896 VSS.n834 53.3664
R5870 VSS.n4900 VSS.n835 53.3664
R5871 VSS.n4869 VSS.n4868 53.3664
R5872 VSS.n1001 VSS.n989 53.3664
R5873 VSS.n4855 VSS.n988 53.3664
R5874 VSS.n3719 VSS.n987 53.3664
R5875 VSS.n3699 VSS.n982 53.3664
R5876 VSS.n3695 VSS.n983 53.3664
R5877 VSS.n3691 VSS.n984 53.3664
R5878 VSS.n3687 VSS.n985 53.3664
R5879 VSS.n4883 VSS.n841 53.3664
R5880 VSS.n4870 VSS.n979 53.3664
R5881 VSS.n980 VSS.n977 53.3664
R5882 VSS.n3471 VSS.n981 53.3664
R5883 VSS.n4808 VSS.n990 53.3664
R5884 VSS.n4807 VSS.n991 53.3664
R5885 VSS.n4803 VSS.n992 53.3664
R5886 VSS.n4799 VSS.n993 53.3664
R5887 VSS.n995 VSS.n990 53.3664
R5888 VSS.n4804 VSS.n991 53.3664
R5889 VSS.n4800 VSS.n992 53.3664
R5890 VSS.n4796 VSS.n993 53.3664
R5891 VSS.n4888 VSS.n832 53.3664
R5892 VSS.n4895 VSS.n833 53.3664
R5893 VSS.n4899 VSS.n834 53.3664
R5894 VSS.n4902 VSS.n835 53.3664
R5895 VSS.n3452 VSS.n821 53.3664
R5896 VSS.n3461 VSS.n828 53.3664
R5897 VSS.n4875 VSS.n820 53.3664
R5898 VSS.n843 VSS.n831 53.3664
R5899 VSS.n3686 VSS.n981 53.3664
R5900 VSS.n3470 VSS.n980 53.3664
R5901 VSS.n4871 VSS.n4870 53.3664
R5902 VSS.n978 VSS.n841 53.3664
R5903 VSS.n1030 VSS.n1014 53.3664
R5904 VSS.n3781 VSS.n1015 53.3664
R5905 VSS.n3789 VSS.n1016 53.3664
R5906 VSS.n3797 VSS.n1018 53.3664
R5907 VSS.n4826 VSS.n1025 53.3664
R5908 VSS.n4825 VSS.n1026 53.3664
R5909 VSS.n4821 VSS.n1027 53.3664
R5910 VSS.n4817 VSS.n1028 53.3664
R5911 VSS.n1029 VSS.n1025 53.3664
R5912 VSS.n4822 VSS.n1026 53.3664
R5913 VSS.n4818 VSS.n1027 53.3664
R5914 VSS.n4814 VSS.n1028 53.3664
R5915 VSS.n4864 VSS.n999 53.3664
R5916 VSS.n4851 VSS.n1013 53.3664
R5917 VSS.n1017 VSS.n1011 53.3664
R5918 VSS.n3751 VSS.n1021 53.3664
R5919 VSS.n3747 VSS.n1022 53.3664
R5920 VSS.n3743 VSS.n1023 53.3664
R5921 VSS.n3739 VSS.n1024 53.3664
R5922 VSS.n3742 VSS.n1024 53.3664
R5923 VSS.n3746 VSS.n1023 53.3664
R5924 VSS.n3750 VSS.n1022 53.3664
R5925 VSS.n3802 VSS.n1021 53.3664
R5926 VSS.n3690 VSS.n985 53.3664
R5927 VSS.n3694 VSS.n984 53.3664
R5928 VSS.n3698 VSS.n983 53.3664
R5929 VSS.n3702 VSS.n982 53.3664
R5930 VSS.n3727 VSS.n987 53.3664
R5931 VSS.n3718 VSS.n988 53.3664
R5932 VSS.n4856 VSS.n989 53.3664
R5933 VSS.n4869 VSS.n994 53.3664
R5934 VSS.n3709 VSS.n1017 53.3664
R5935 VSS.n4852 VSS.n4851 53.3664
R5936 VSS.n1012 VSS.n999 53.3664
R5937 VSS.n932 VSS.n449 53.3664
R5938 VSS.n923 VSS.n450 53.3664
R5939 VSS.n5109 VSS.n451 53.3664
R5940 VSS.n5122 VSS.n456 53.3664
R5941 VSS.n914 VSS.n476 53.3664
R5942 VSS.n5105 VSS.n5104 53.3664
R5943 VSS.n471 VSS.n461 53.3664
R5944 VSS.n2078 VSS.n259 53.3664
R5945 VSS.n2236 VSS.n247 53.3664
R5946 VSS.n2089 VSS.n256 53.3664
R5947 VSS.n2222 VSS.n248 53.3664
R5948 VSS.n5305 VSS.n5304 53.3664
R5949 VSS.n264 VSS.n262 53.3664
R5950 VSS.n5299 VSS.n261 53.3664
R5951 VSS.n5295 VSS.n260 53.3664
R5952 VSS.n5305 VSS.n263 53.3664
R5953 VSS.n5300 VSS.n262 53.3664
R5954 VSS.n5296 VSS.n261 53.3664
R5955 VSS.n5292 VSS.n260 53.3664
R5956 VSS.n258 VSS.n244 53.3664
R5957 VSS.n5273 VSS.n257 53.3664
R5958 VSS.n286 VSS.n255 53.3664
R5959 VSS.n2202 VSS.n253 53.3664
R5960 VSS.n2198 VSS.n252 53.3664
R5961 VSS.n2194 VSS.n251 53.3664
R5962 VSS.n2190 VSS.n250 53.3664
R5963 VSS.n2739 VSS.n2738 53.3664
R5964 VSS.n2141 VSS.n2071 53.3664
R5965 VSS.n2144 VSS.n2143 53.3664
R5966 VSS.n2167 VSS.n2166 53.3664
R5967 VSS.n2735 VSS.n2734 53.3664
R5968 VSS.n2729 VSS.n2073 53.3664
R5969 VSS.n2728 VSS.n2727 53.3664
R5970 VSS.n2721 VSS.n2075 53.3664
R5971 VSS.n2736 VSS.n2735 53.3664
R5972 VSS.n2730 VSS.n2729 53.3664
R5973 VSS.n2727 VSS.n2726 53.3664
R5974 VSS.n2722 VSS.n2721 53.3664
R5975 VSS.n2232 VSS.n2077 53.3664
R5976 VSS.n2231 VSS.n2086 53.3664
R5977 VSS.n2218 VSS.n2217 53.3664
R5978 VSS.n2169 VSS.n2103 53.3664
R5979 VSS.n2176 VSS.n2175 53.3664
R5980 VSS.n2177 VSS.n2101 53.3664
R5981 VSS.n2184 VSS.n2183 53.3664
R5982 VSS.n2183 VSS.n2182 53.3664
R5983 VSS.n2178 VSS.n2177 53.3664
R5984 VSS.n2175 VSS.n2174 53.3664
R5985 VSS.n2170 VSS.n2169 53.3664
R5986 VSS.n2193 VSS.n250 53.3664
R5987 VSS.n2197 VSS.n251 53.3664
R5988 VSS.n2201 VSS.n252 53.3664
R5989 VSS.n2204 VSS.n253 53.3664
R5990 VSS.n2855 VSS.n508 53.3664
R5991 VSS.n3014 VSS.n496 53.3664
R5992 VSS.n2866 VSS.n505 53.3664
R5993 VSS.n3000 VSS.n497 53.3664
R5994 VSS.n5098 VSS.n5097 53.3664
R5995 VSS.n513 VSS.n511 53.3664
R5996 VSS.n5092 VSS.n510 53.3664
R5997 VSS.n5088 VSS.n509 53.3664
R5998 VSS.n5098 VSS.n512 53.3664
R5999 VSS.n5093 VSS.n511 53.3664
R6000 VSS.n5089 VSS.n510 53.3664
R6001 VSS.n5085 VSS.n509 53.3664
R6002 VSS.n507 VSS.n493 53.3664
R6003 VSS.n5066 VSS.n506 53.3664
R6004 VSS.n714 VSS.n504 53.3664
R6005 VSS.n2981 VSS.n502 53.3664
R6006 VSS.n2977 VSS.n501 53.3664
R6007 VSS.n2973 VSS.n500 53.3664
R6008 VSS.n2969 VSS.n499 53.3664
R6009 VSS.n3045 VSS.n3044 53.3664
R6010 VSS.n2920 VSS.n2028 53.3664
R6011 VSS.n2923 VSS.n2922 53.3664
R6012 VSS.n2946 VSS.n2945 53.3664
R6013 VSS.n3041 VSS.n3040 53.3664
R6014 VSS.n3035 VSS.n2850 53.3664
R6015 VSS.n3034 VSS.n3033 53.3664
R6016 VSS.n3027 VSS.n2852 53.3664
R6017 VSS.n3042 VSS.n3041 53.3664
R6018 VSS.n3036 VSS.n3035 53.3664
R6019 VSS.n3033 VSS.n3032 53.3664
R6020 VSS.n3028 VSS.n3027 53.3664
R6021 VSS.n3010 VSS.n2854 53.3664
R6022 VSS.n3009 VSS.n2863 53.3664
R6023 VSS.n2996 VSS.n2995 53.3664
R6024 VSS.n2948 VSS.n2882 53.3664
R6025 VSS.n2955 VSS.n2954 53.3664
R6026 VSS.n2956 VSS.n2880 53.3664
R6027 VSS.n2963 VSS.n2962 53.3664
R6028 VSS.n2962 VSS.n2961 53.3664
R6029 VSS.n2957 VSS.n2956 53.3664
R6030 VSS.n2954 VSS.n2953 53.3664
R6031 VSS.n2949 VSS.n2948 53.3664
R6032 VSS.n2972 VSS.n499 53.3664
R6033 VSS.n2976 VSS.n500 53.3664
R6034 VSS.n2980 VSS.n501 53.3664
R6035 VSS.n2983 VSS.n502 53.3664
R6036 VSS.n2875 VSS.n497 53.3664
R6037 VSS.n3001 VSS.n505 53.3664
R6038 VSS.n2865 VSS.n496 53.3664
R6039 VSS.n3015 VSS.n508 53.3664
R6040 VSS.n2997 VSS.n2996 53.3664
R6041 VSS.n2994 VSS.n2863 53.3664
R6042 VSS.n3011 VSS.n3010 53.3664
R6043 VSS.n2098 VSS.n248 53.3664
R6044 VSS.n2223 VSS.n256 53.3664
R6045 VSS.n2088 VSS.n247 53.3664
R6046 VSS.n2237 VSS.n259 53.3664
R6047 VSS.n2219 VSS.n2218 53.3664
R6048 VSS.n2216 VSS.n2086 53.3664
R6049 VSS.n2233 VSS.n2232 53.3664
R6050 VSS.n3278 VSS.n1528 53.3664
R6051 VSS.n3411 VSS.n1516 53.3664
R6052 VSS.n3289 VSS.n1525 53.3664
R6053 VSS.n3397 VSS.n1517 53.3664
R6054 VSS.n4472 VSS.n4471 53.3664
R6055 VSS.n1533 VSS.n1531 53.3664
R6056 VSS.n4466 VSS.n1530 53.3664
R6057 VSS.n4462 VSS.n1529 53.3664
R6058 VSS.n4472 VSS.n1532 53.3664
R6059 VSS.n4467 VSS.n1531 53.3664
R6060 VSS.n4463 VSS.n1530 53.3664
R6061 VSS.n4459 VSS.n1529 53.3664
R6062 VSS.n1527 VSS.n1513 53.3664
R6063 VSS.n4440 VSS.n1526 53.3664
R6064 VSS.n1551 VSS.n1524 53.3664
R6065 VSS.n3378 VSS.n1522 53.3664
R6066 VSS.n3374 VSS.n1521 53.3664
R6067 VSS.n3370 VSS.n1520 53.3664
R6068 VSS.n3366 VSS.n1519 53.3664
R6069 VSS.n3953 VSS.n3952 53.3664
R6070 VSS.n3323 VSS.n1952 53.3664
R6071 VSS.n3326 VSS.n3325 53.3664
R6072 VSS.n3343 VSS.n3342 53.3664
R6073 VSS.n3949 VSS.n3948 53.3664
R6074 VSS.n3943 VSS.n3273 53.3664
R6075 VSS.n3942 VSS.n3941 53.3664
R6076 VSS.n3935 VSS.n3275 53.3664
R6077 VSS.n3950 VSS.n3949 53.3664
R6078 VSS.n3944 VSS.n3943 53.3664
R6079 VSS.n3941 VSS.n3940 53.3664
R6080 VSS.n3936 VSS.n3935 53.3664
R6081 VSS.n3407 VSS.n3277 53.3664
R6082 VSS.n3406 VSS.n3286 53.3664
R6083 VSS.n3393 VSS.n3392 53.3664
R6084 VSS.n3345 VSS.n3305 53.3664
R6085 VSS.n3352 VSS.n3351 53.3664
R6086 VSS.n3353 VSS.n3303 53.3664
R6087 VSS.n3360 VSS.n3359 53.3664
R6088 VSS.n3359 VSS.n3358 53.3664
R6089 VSS.n3354 VSS.n3353 53.3664
R6090 VSS.n3351 VSS.n3350 53.3664
R6091 VSS.n3346 VSS.n3345 53.3664
R6092 VSS.n3369 VSS.n1519 53.3664
R6093 VSS.n3373 VSS.n1520 53.3664
R6094 VSS.n3377 VSS.n1521 53.3664
R6095 VSS.n3380 VSS.n1522 53.3664
R6096 VSS.n3298 VSS.n1517 53.3664
R6097 VSS.n3398 VSS.n1525 53.3664
R6098 VSS.n3288 VSS.n1516 53.3664
R6099 VSS.n3412 VSS.n1528 53.3664
R6100 VSS.n3394 VSS.n3393 53.3664
R6101 VSS.n3391 VSS.n3286 53.3664
R6102 VSS.n3408 VSS.n3407 53.3664
R6103 VSS.n3857 VSS.n1038 53.3664
R6104 VSS.n3849 VSS.n1046 53.3664
R6105 VSS.n3840 VSS.n1037 53.3664
R6106 VSS.n4785 VSS.n1049 53.3664
R6107 VSS.n3832 VSS.n1072 53.3664
R6108 VSS.n3837 VSS.n1070 53.3664
R6109 VSS.n4781 VSS.n4780 53.3664
R6110 VSS.n2657 VSS.n2058 53.3664
R6111 VSS.n2631 VSS.n2047 53.3664
R6112 VSS.n2646 VSS.n2055 53.3664
R6113 VSS.n2637 VSS.n2048 53.3664
R6114 VSS.n2106 VSS.n2052 53.3664
R6115 VSS.n2110 VSS.n2051 53.3664
R6116 VSS.n2114 VSS.n2050 53.3664
R6117 VSS.n2118 VSS.n2049 53.3664
R6118 VSS.n2115 VSS.n2049 53.3664
R6119 VSS.n2111 VSS.n2050 53.3664
R6120 VSS.n2107 VSS.n2051 53.3664
R6121 VSS.n2052 VSS.n2045 53.3664
R6122 VSS.n2069 VSS.n2057 53.3664
R6123 VSS.n2138 VSS.n2056 53.3664
R6124 VSS.n2148 VSS.n2054 53.3664
R6125 VSS.n2661 VSS.n2059 53.3664
R6126 VSS.n2662 VSS.n2060 53.3664
R6127 VSS.n2666 VSS.n2061 53.3664
R6128 VSS.n2670 VSS.n2062 53.3664
R6129 VSS.n2658 VSS.n2059 53.3664
R6130 VSS.n2665 VSS.n2060 53.3664
R6131 VSS.n2669 VSS.n2061 53.3664
R6132 VSS.n2672 VSS.n2062 53.3664
R6133 VSS.n2048 VSS.n2044 53.3664
R6134 VSS.n2636 VSS.n2055 53.3664
R6135 VSS.n2647 VSS.n2047 53.3664
R6136 VSS.n2630 VSS.n2058 53.3664
R6137 VSS.n2005 VSS.n2001 53.3664
R6138 VSS.n2805 VSS.n2012 53.3664
R6139 VSS.n2816 VSS.n2004 53.3664
R6140 VSS.n2799 VSS.n2015 53.3664
R6141 VSS.n3140 VSS.n1095 53.3664
R6142 VSS.n3136 VSS.n1103 53.3664
R6143 VSS.n3125 VSS.n1094 53.3664
R6144 VSS.n3120 VSS.n1106 53.3664
R6145 VSS.n3228 VSS.n1929 53.3664
R6146 VSS.n3200 VSS.n1936 53.3664
R6147 VSS.n3239 VSS.n1928 53.3664
R6148 VSS.n3191 VSS.n1939 53.3664
R6149 VSS.n4126 VSS.n1815 53.3664
R6150 VSS.n4116 VSS.n1823 53.3664
R6151 VSS.n4111 VSS.n1814 53.3664
R6152 VSS.n4100 VSS.n1826 53.3664
R6153 VSS.n2168 VSS.n2167 53.3664
R6154 VSS.n2143 VSS.n2123 53.3664
R6155 VSS.n2142 VSS.n2141 53.3664
R6156 VSS.n2740 VSS.n2739 53.3664
R6157 VSS.n2947 VSS.n2946 53.3664
R6158 VSS.n2922 VSS.n2902 53.3664
R6159 VSS.n2921 VSS.n2920 53.3664
R6160 VSS.n3046 VSS.n3045 53.3664
R6161 VSS.n3414 VSS.n1073 53.3664
R6162 VSS.n4744 VSS.n1071 53.3664
R6163 VSS.n1143 VSS.n1069 53.3664
R6164 VSS.n4757 VSS.n1068 53.3664
R6165 VSS.n3344 VSS.n3343 53.3664
R6166 VSS.n3325 VSS.n3306 53.3664
R6167 VSS.n3324 VSS.n3323 53.3664
R6168 VSS.n3954 VSS.n3953 53.3664
R6169 VSS.n1845 VSS.n1793 53.3664
R6170 VSS.n4231 VSS.n1801 53.3664
R6171 VSS.n4243 VSS.n1792 53.3664
R6172 VSS.n2163 VSS.n2054 53.3664
R6173 VSS.n2147 VSS.n2056 53.3664
R6174 VSS.n2137 VSS.n2057 53.3664
R6175 VSS.n2942 VSS.n2011 53.3664
R6176 VSS.n2926 VSS.n2013 53.3664
R6177 VSS.n2916 VSS.n2014 53.3664
R6178 VSS.n4740 VSS.n1102 53.3664
R6179 VSS.n1147 VSS.n1104 53.3664
R6180 VSS.n4753 VSS.n1105 53.3664
R6181 VSS.n1935 VSS.n1925 53.3664
R6182 VSS.n3329 VSS.n1937 53.3664
R6183 VSS.n3319 VSS.n1938 53.3664
R6184 VSS.n4218 VSS.n1822 53.3664
R6185 VSS.n4227 VSS.n1824 53.3664
R6186 VSS.n4239 VSS.n1825 53.3664
R6187 VSS.n4267 VSS.n1804 53.3664
R6188 VSS.n4263 VSS.n1805 53.3664
R6189 VSS.n4259 VSS.n1806 53.3664
R6190 VSS.n4281 VSS.n1807 53.3664
R6191 VSS.n4337 VSS.n1777 53.3664
R6192 VSS.n4332 VSS.n1776 53.3664
R6193 VSS.n4328 VSS.n1775 53.3664
R6194 VSS.n4324 VSS.n1774 53.3664
R6195 VSS.n2480 VSS.n1765 53.3664
R6196 VSS.n2471 VSS.n1772 53.3664
R6197 VSS.n2462 VSS.n1763 53.3664
R6198 VSS.n4289 VSS.n1773 53.3664
R6199 VSS.n2486 VSS.n1800 53.3664
R6200 VSS.n2456 VSS.n1802 53.3664
R6201 VSS.n4284 VSS.n1791 53.3664
R6202 VSS.n4283 VSS.n1790 53.3664
R6203 VSS.n2505 VSS.n1771 53.3664
R6204 VSS.n2501 VSS.n1770 53.3664
R6205 VSS.n2497 VSS.n1769 53.3664
R6206 VSS.n2493 VSS.n1768 53.3664
R6207 VSS.n2394 VSS.n1740 53.3664
R6208 VSS.n2398 VSS.n1710 53.3664
R6209 VSS.n2402 VSS.n1709 53.3664
R6210 VSS.n2406 VSS.n1708 53.3664
R6211 VSS.n532 VSS.n228 53.3664
R6212 VSS.n5265 VSS.n227 53.3664
R6213 VSS.n281 VSS.n222 53.3664
R6214 VSS.n5278 VSS.n221 53.3664
R6215 VSS.n891 VSS.n477 53.3664
R6216 VSS.n5058 VSS.n475 53.3664
R6217 VSS.n709 VSS.n474 53.3664
R6218 VSS.n5071 VSS.n473 53.3664
R6219 VSS.n3803 VSS.n1018 53.3664
R6220 VSS.n3796 VSS.n1016 53.3664
R6221 VSS.n3788 VSS.n1015 53.3664
R6222 VSS.n3780 VSS.n1014 53.3664
R6223 VSS.n1585 VSS.n1497 53.3664
R6224 VSS.n4432 VSS.n1495 53.3664
R6225 VSS.n1546 VSS.n1494 53.3664
R6226 VSS.n4445 VSS.n1493 53.3664
R6227 VSS.n2432 VSS.n1742 53.3664
R6228 VSS.n2424 VSS.n1743 53.3664
R6229 VSS.n4345 VSS.n1744 53.3664
R6230 VSS.n4361 VSS.n1749 53.3664
R6231 VSS.n5261 VSS.n255 53.3664
R6232 VSS.n285 VSS.n257 53.3664
R6233 VSS.n5274 VSS.n258 53.3664
R6234 VSS.n5054 VSS.n504 53.3664
R6235 VSS.n713 VSS.n506 53.3664
R6236 VSS.n5067 VSS.n507 53.3664
R6237 VSS.n3800 VSS.n1045 53.3664
R6238 VSS.n3792 VSS.n1047 53.3664
R6239 VSS.n3784 VSS.n1048 53.3664
R6240 VSS.n4428 VSS.n1524 53.3664
R6241 VSS.n1550 VSS.n1526 53.3664
R6242 VSS.n4441 VSS.n1527 53.3664
R6243 VSS.n2509 VSS.n1766 53.3664
R6244 VSS.n2428 VSS.n1764 53.3664
R6245 VSS.n4342 VSS.n4341 53.3664
R6246 VSS.n4339 VSS.n1754 53.3664
R6247 VSS.n113 VSS.n103 53.3664
R6248 VSS.n5390 VSS.n115 53.3664
R6249 VSS.n5403 VSS.n116 53.3664
R6250 VSS.n412 VSS.n402 53.3664
R6251 VSS.n5177 VSS.n414 53.3664
R6252 VSS.n5190 VSS.n415 53.3664
R6253 VSS.n827 VSS.n817 53.3664
R6254 VSS.n4924 VSS.n829 53.3664
R6255 VSS.n4937 VSS.n830 53.3664
R6256 VSS.n3648 VSS.n3514 53.3664
R6257 VSS.n3641 VSS.n3563 53.3664
R6258 VSS.n3659 VSS.n3564 53.3664
R6259 VSS.n5504 VSS.n5503 53.3664
R6260 VSS.n5501 VSS.n5500 53.3664
R6261 VSS.n5484 VSS.n46 53.3664
R6262 VSS.n4628 VSS.t88 52.4309
R6263 VSS.n4624 VSS.t15 52.242
R6264 VSS.n323 VSS.n320 49.7381
R6265 VSS.n330 VSS.n324 49.7381
R6266 VSS.n764 VSS.n325 49.7381
R6267 VSS.n1653 VSS.n326 49.7381
R6268 VSS.n81 VSS.n75 49.7381
R6269 VSS.n5217 VSS.n76 49.7381
R6270 VSS.n4964 VSS.n77 49.7381
R6271 VSS.n5438 VSS.n5437 49.7381
R6272 VSS.n698 VSS.n300 49.7381
R6273 VSS.n5012 VSS.n728 49.7381
R6274 VSS.n736 VSS.n732 49.7381
R6275 VSS.n1564 VSS.n733 49.7381
R6276 VSS.n4689 VSS.n4688 49.7381
R6277 VSS.n1305 VSS.n1304 49.7381
R6278 VSS.n3919 VSS.n3904 49.7381
R6279 VSS.n4049 VSS.n4009 49.7381
R6280 VSS.n1202 VSS.n1198 49.7381
R6281 VSS.n1193 VSS.n1130 49.7381
R6282 VSS.n1166 VSS.n1165 49.7381
R6283 VSS.n3973 VSS.n1199 49.7381
R6284 VSS.n5235 VSS.n323 48.7629
R6285 VSS.n5233 VSS.n330 48.7629
R6286 VSS.n764 VSS.n328 48.7629
R6287 VSS.n1653 VSS.n327 48.7629
R6288 VSS.n5435 VSS.n81 48.7629
R6289 VSS.n5217 VSS.n79 48.7629
R6290 VSS.n4964 VSS.n78 48.7629
R6291 VSS.n5438 VSS.n72 48.7629
R6292 VSS.n300 VSS.n296 48.7629
R6293 VSS.n728 VSS.n724 48.7629
R6294 VSS.n5010 VSS.n736 48.7629
R6295 VSS.n1564 VSS.n734 48.7629
R6296 VSS.n4689 VSS.n1221 48.7629
R6297 VSS.n1305 VSS.n1276 48.7629
R6298 VSS.n3921 VSS.n3904 48.7629
R6299 VSS.n4050 VSS.n4049 48.7629
R6300 VSS.n4712 VSS.n1202 48.7629
R6301 VSS.n4714 VSS.n1193 48.7629
R6302 VSS.n1166 VSS.n1158 48.7629
R6303 VSS.n3973 VSS.n1200 48.7629
R6304 VSS.n1376 VSS.t10 42.6154
R6305 VSS.n1398 VSS.t18 42.5516
R6306 VSS.n1375 VSS.t9 42.4377
R6307 VSS.n4622 VSS.t17 42.3691
R6308 VSS.n1565 VSS.n1561 40.8246
R6309 VSS.n4417 VSS.n4416 40.8246
R6310 VSS.n4413 VSS.n1572 40.8246
R6311 VSS.n4411 VSS.n1571 40.8246
R6312 VSS.n4410 VSS.n4409 40.8246
R6313 VSS.n1576 VSS.n1570 40.8246
R6314 VSS.n1578 VSS.n1574 40.8246
R6315 VSS.n1580 VSS.n1569 40.8246
R6316 VSS.n1582 VSS.n1575 40.8246
R6317 VSS.n4406 VSS.n1568 40.8246
R6318 VSS.n4407 VSS.n1567 40.8246
R6319 VSS.n301 VSS.n297 40.8246
R6320 VSS.n5250 VSS.n5249 40.8246
R6321 VSS.n5246 VSS.n308 40.8246
R6322 VSS.n5244 VSS.n307 40.8246
R6323 VSS.n5243 VSS.n5242 40.8246
R6324 VSS.n312 VSS.n306 40.8246
R6325 VSS.n314 VSS.n310 40.8246
R6326 VSS.n316 VSS.n305 40.8246
R6327 VSS.n318 VSS.n311 40.8246
R6328 VSS.n5239 VSS.n304 40.8246
R6329 VSS.n5240 VSS.n303 40.8246
R6330 VSS.n5226 VSS.n336 40.8246
R6331 VSS.n5226 VSS.n5225 40.8246
R6332 VSS.n347 VSS.n344 40.8246
R6333 VSS.n347 VSS.n339 40.8246
R6334 VSS.n351 VSS.n345 40.8246
R6335 VSS.n351 VSS.n340 40.8246
R6336 VSS.n357 VSS.n356 40.8246
R6337 VSS.n356 VSS.n341 40.8246
R6338 VSS.n5222 VSS.n5221 40.8246
R6339 VSS.n5218 VSS.n338 40.8246
R6340 VSS.n336 VSS.n334 40.8246
R6341 VSS.n5221 VSS.n338 40.8246
R6342 VSS.n5223 VSS.n5222 40.8246
R6343 VSS.n342 VSS.n341 40.8246
R6344 VSS.n346 VSS.n340 40.8246
R6345 VSS.n357 VSS.n346 40.8246
R6346 VSS.n349 VSS.n339 40.8246
R6347 VSS.n349 VSS.n345 40.8246
R6348 VSS.n5225 VSS.n337 40.8246
R6349 VSS.n344 VSS.n337 40.8246
R6350 VSS.n5216 VSS.n360 40.8246
R6351 VSS.n376 VSS.n362 40.8246
R6352 VSS.n376 VSS.n371 40.8246
R6353 VSS.n380 VSS.n363 40.8246
R6354 VSS.n380 VSS.n372 40.8246
R6355 VSS.n373 VSS.n364 40.8246
R6356 VSS.n387 VSS.n373 40.8246
R6357 VSS.n370 VSS.n365 40.8246
R6358 VSS.n389 VSS.n370 40.8246
R6359 VSS.n392 VSS.n366 40.8246
R6360 VSS.n5214 VSS.n367 40.8246
R6361 VSS.n5212 VSS.n368 40.8246
R6362 VSS.n392 VSS.n367 40.8246
R6363 VSS.n390 VSS.n389 40.8246
R6364 VSS.n390 VSS.n366 40.8246
R6365 VSS.n387 VSS.n386 40.8246
R6366 VSS.n386 VSS.n365 40.8246
R6367 VSS.n382 VSS.n372 40.8246
R6368 VSS.n382 VSS.n364 40.8246
R6369 VSS.n378 VSS.n371 40.8246
R6370 VSS.n378 VSS.n363 40.8246
R6371 VSS.n374 VSS.n360 40.8246
R6372 VSS.n374 VSS.n362 40.8246
R6373 VSS.n4963 VSS.n775 40.8246
R6374 VSS.n791 VSS.n777 40.8246
R6375 VSS.n791 VSS.n786 40.8246
R6376 VSS.n795 VSS.n778 40.8246
R6377 VSS.n795 VSS.n787 40.8246
R6378 VSS.n788 VSS.n779 40.8246
R6379 VSS.n802 VSS.n788 40.8246
R6380 VSS.n785 VSS.n780 40.8246
R6381 VSS.n804 VSS.n785 40.8246
R6382 VSS.n807 VSS.n781 40.8246
R6383 VSS.n4961 VSS.n782 40.8246
R6384 VSS.n4959 VSS.n783 40.8246
R6385 VSS.n807 VSS.n782 40.8246
R6386 VSS.n805 VSS.n804 40.8246
R6387 VSS.n805 VSS.n781 40.8246
R6388 VSS.n802 VSS.n801 40.8246
R6389 VSS.n801 VSS.n780 40.8246
R6390 VSS.n797 VSS.n787 40.8246
R6391 VSS.n797 VSS.n779 40.8246
R6392 VSS.n793 VSS.n786 40.8246
R6393 VSS.n793 VSS.n778 40.8246
R6394 VSS.n789 VSS.n775 40.8246
R6395 VSS.n789 VSS.n777 40.8246
R6396 VSS.n741 VSS.n738 40.8246
R6397 VSS.n5006 VSS.n5005 40.8246
R6398 VSS.n5002 VSS.n748 40.8246
R6399 VSS.n5000 VSS.n747 40.8246
R6400 VSS.n4999 VSS.n4998 40.8246
R6401 VSS.n752 VSS.n746 40.8246
R6402 VSS.n754 VSS.n750 40.8246
R6403 VSS.n756 VSS.n745 40.8246
R6404 VSS.n758 VSS.n751 40.8246
R6405 VSS.n4995 VSS.n744 40.8246
R6406 VSS.n4996 VSS.n743 40.8246
R6407 VSS.n2362 VSS.n2361 40.8246
R6408 VSS.n2360 VSS.n2359 40.8246
R6409 VSS.n5323 VSS.n208 40.8246
R6410 VSS.n5322 VSS.n5321 40.8246
R6411 VSS.n5320 VSS.n5319 40.8246
R6412 VSS.n617 VSS.n212 40.8246
R6413 VSS.n619 VSS.n618 40.8246
R6414 VSS.n621 VSS.n620 40.8246
R6415 VSS.n633 VSS.n615 40.8246
R6416 VSS.n636 VSS.n634 40.8246
R6417 VSS.n636 VSS.n635 40.8246
R6418 VSS.n642 VSS.n641 40.8246
R6419 VSS.n640 VSS.n639 40.8246
R6420 VSS.n5114 VSS.n465 40.8246
R6421 VSS.n5113 VSS.n5112 40.8246
R6422 VSS.n918 VSS.n466 40.8246
R6423 VSS.n920 VSS.n919 40.8246
R6424 VSS.n927 VSS.n916 40.8246
R6425 VSS.n929 VSS.n928 40.8246
R6426 VSS.n936 VSS.n912 40.8246
R6427 VSS.n939 VSS.n937 40.8246
R6428 VSS.n938 VSS.n329 40.8246
R6429 VSS.n1003 VSS.n333 40.8246
R6430 VSS.n1005 VSS.n1004 40.8246
R6431 VSS.n4861 VSS.n1006 40.8246
R6432 VSS.n4860 VSS.n4859 40.8246
R6433 VSS.n3713 VSS.n1007 40.8246
R6434 VSS.n3715 VSS.n3714 40.8246
R6435 VSS.n3722 VSS.n3711 40.8246
R6436 VSS.n3724 VSS.n3723 40.8246
R6437 VSS.n3731 VSS.n3707 40.8246
R6438 VSS.n3734 VSS.n3732 40.8246
R6439 VSS.n3733 VSS.n760 40.8246
R6440 VSS.n1482 VSS.n762 40.8246
R6441 VSS.n1484 VSS.n1483 40.8246
R6442 VSS.n4488 VSS.n1485 40.8246
R6443 VSS.n4487 VSS.n4486 40.8246
R6444 VSS.n1627 VSS.n1486 40.8246
R6445 VSS.n1629 VSS.n1628 40.8246
R6446 VSS.n1636 VSS.n1625 40.8246
R6447 VSS.n1638 VSS.n1637 40.8246
R6448 VSS.n1645 VSS.n1621 40.8246
R6449 VSS.n1648 VSS.n1646 40.8246
R6450 VSS.n1647 VSS.n1584 40.8246
R6451 VSS.n4400 VSS.n4399 40.8246
R6452 VSS.n1697 VSS.n1688 40.8246
R6453 VSS.n4374 VSS.n1698 40.8246
R6454 VSS.n4373 VSS.n4372 40.8246
R6455 VSS.n4371 VSS.n4370 40.8246
R6456 VSS.n1716 VSS.n1700 40.8246
R6457 VSS.n1715 VSS.n1714 40.8246
R6458 VSS.n1729 VSS.n1712 40.8246
R6459 VSS.n1734 VSS.n1730 40.8246
R6460 VSS.n1733 VSS.n1732 40.8246
R6461 VSS.n1732 VSS.n1731 40.8246
R6462 VSS.n2361 VSS.n2360 40.8246
R6463 VSS.n5323 VSS.n5322 40.8246
R6464 VSS.n5319 VSS.n212 40.8246
R6465 VSS.n620 VSS.n619 40.8246
R6466 VSS.n634 VSS.n633 40.8246
R6467 VSS.n639 VSS.n465 40.8246
R6468 VSS.n5112 VSS.n466 40.8246
R6469 VSS.n920 VSS.n916 40.8246
R6470 VSS.n929 VSS.n912 40.8246
R6471 VSS.n939 VSS.n938 40.8246
R6472 VSS.n5230 VSS.n333 40.8246
R6473 VSS.n1006 VSS.n1005 40.8246
R6474 VSS.n4859 VSS.n1007 40.8246
R6475 VSS.n3715 VSS.n3711 40.8246
R6476 VSS.n3724 VSS.n3707 40.8246
R6477 VSS.n3734 VSS.n3733 40.8246
R6478 VSS.n4990 VSS.n762 40.8246
R6479 VSS.n1485 VSS.n1484 40.8246
R6480 VSS.n4486 VSS.n1486 40.8246
R6481 VSS.n1629 VSS.n1625 40.8246
R6482 VSS.n1638 VSS.n1621 40.8246
R6483 VSS.n1648 VSS.n1647 40.8246
R6484 VSS.n4399 VSS.n1688 40.8246
R6485 VSS.n4374 VSS.n4373 40.8246
R6486 VSS.n4370 VSS.n1700 40.8246
R6487 VSS.n1714 VSS.n1712 40.8246
R6488 VSS.n1734 VSS.n1733 40.8246
R6489 VSS.n1730 VSS.n1729 40.8246
R6490 VSS.n1716 VSS.n1715 40.8246
R6491 VSS.n4372 VSS.n4371 40.8246
R6492 VSS.n1698 VSS.n1697 40.8246
R6493 VSS.n4401 VSS.n4400 40.8246
R6494 VSS.n1646 VSS.n1645 40.8246
R6495 VSS.n1637 VSS.n1636 40.8246
R6496 VSS.n1628 VSS.n1627 40.8246
R6497 VSS.n4488 VSS.n4487 40.8246
R6498 VSS.n1483 VSS.n1482 40.8246
R6499 VSS.n3732 VSS.n3731 40.8246
R6500 VSS.n3723 VSS.n3722 40.8246
R6501 VSS.n3714 VSS.n3713 40.8246
R6502 VSS.n4861 VSS.n4860 40.8246
R6503 VSS.n1004 VSS.n1003 40.8246
R6504 VSS.n937 VSS.n936 40.8246
R6505 VSS.n928 VSS.n927 40.8246
R6506 VSS.n919 VSS.n918 40.8246
R6507 VSS.n5114 VSS.n5113 40.8246
R6508 VSS.n641 VSS.n640 40.8246
R6509 VSS.n621 VSS.n615 40.8246
R6510 VSS.n618 VSS.n617 40.8246
R6511 VSS.n5321 VSS.n5320 40.8246
R6512 VSS.n2359 VSS.n208 40.8246
R6513 VSS.n2363 VSS.n2362 40.8246
R6514 VSS.n5442 VSS.n65 40.8246
R6515 VSS.n5444 VSS.n5443 40.8246
R6516 VSS.n5447 VSS.n66 40.8246
R6517 VSS.n5449 VSS.n5448 40.8246
R6518 VSS.n5452 VSS.n67 40.8246
R6519 VSS.n5454 VSS.n5453 40.8246
R6520 VSS.n5456 VSS.n68 40.8246
R6521 VSS.n5459 VSS.n69 40.8246
R6522 VSS.n5461 VSS.n5460 40.8246
R6523 VSS.n5465 VSS.n64 40.8246
R6524 VSS.n5464 VSS.n5463 40.8246
R6525 VSS.n5473 VSS.n59 40.8246
R6526 VSS.n2283 VSS.n2282 40.8246
R6527 VSS.n2281 VSS.n2280 40.8246
R6528 VSS.n5343 VSS.n177 40.8246
R6529 VSS.n5342 VSS.n5341 40.8246
R6530 VSS.n5340 VSS.n5339 40.8246
R6531 VSS.n574 VSS.n179 40.8246
R6532 VSS.n581 VSS.n572 40.8246
R6533 VSS.n583 VSS.n582 40.8246
R6534 VSS.n590 VSS.n569 40.8246
R6535 VSS.n593 VSS.n591 40.8246
R6536 VSS.n593 VSS.n592 40.8246
R6537 VSS.n431 VSS.n84 40.8246
R6538 VSS.n433 VSS.n432 40.8246
R6539 VSS.n5133 VSS.n434 40.8246
R6540 VSS.n5132 VSS.n5131 40.8246
R6541 VSS.n852 VSS.n435 40.8246
R6542 VSS.n856 VSS.n853 40.8246
R6543 VSS.n855 VSS.n854 40.8246
R6544 VSS.n869 VSS.n850 40.8246
R6545 VSS.n871 VSS.n870 40.8246
R6546 VSS.n963 VSS.n848 40.8246
R6547 VSS.n965 VSS.n964 40.8246
R6548 VSS.n969 VSS.n968 40.8246
R6549 VSS.n971 VSS.n970 40.8246
R6550 VSS.n4880 VSS.n972 40.8246
R6551 VSS.n4879 VSS.n4878 40.8246
R6552 VSS.n3456 VSS.n973 40.8246
R6553 VSS.n3458 VSS.n3457 40.8246
R6554 VSS.n3465 VSS.n3455 40.8246
R6555 VSS.n3467 VSS.n3466 40.8246
R6556 VSS.n3474 VSS.n3451 40.8246
R6557 VSS.n3683 VSS.n3475 40.8246
R6558 VSS.n3682 VSS.n3681 40.8246
R6559 VSS.n3678 VSS.n3677 40.8246
R6560 VSS.n3676 VSS.n3675 40.8246
R6561 VSS.n3524 VSS.n3480 40.8246
R6562 VSS.n3526 VSS.n3525 40.8246
R6563 VSS.n3533 VSS.n3519 40.8246
R6564 VSS.n3554 VSS.n3534 40.8246
R6565 VSS.n3553 VSS.n3552 40.8246
R6566 VSS.n3551 VSS.n3550 40.8246
R6567 VSS.n3544 VSS.n3535 40.8246
R6568 VSS.n3543 VSS.n3542 40.8246
R6569 VSS.n3541 VSS.n3540 40.8246
R6570 VSS.n4504 VSS.n4503 40.8246
R6571 VSS.n4575 VSS.n1446 40.8246
R6572 VSS.n4574 VSS.n4573 40.8246
R6573 VSS.n4531 VSS.n1447 40.8246
R6574 VSS.n4562 VSS.n4532 40.8246
R6575 VSS.n4561 VSS.n4560 40.8246
R6576 VSS.n4559 VSS.n4558 40.8246
R6577 VSS.n4545 VSS.n4534 40.8246
R6578 VSS.n4547 VSS.n4546 40.8246
R6579 VSS.n5533 VSS.n26 40.8246
R6580 VSS.n5534 VSS.n5533 40.8246
R6581 VSS.n2282 VSS.n2281 40.8246
R6582 VSS.n5343 VSS.n5342 40.8246
R6583 VSS.n5339 VSS.n179 40.8246
R6584 VSS.n582 VSS.n581 40.8246
R6585 VSS.n591 VSS.n590 40.8246
R6586 VSS.n434 VSS.n433 40.8246
R6587 VSS.n5131 VSS.n435 40.8246
R6588 VSS.n856 VSS.n855 40.8246
R6589 VSS.n870 VSS.n869 40.8246
R6590 VSS.n964 VSS.n963 40.8246
R6591 VSS.n968 VSS.n967 40.8246
R6592 VSS.n972 VSS.n971 40.8246
R6593 VSS.n4878 VSS.n973 40.8246
R6594 VSS.n3458 VSS.n3455 40.8246
R6595 VSS.n3467 VSS.n3451 40.8246
R6596 VSS.n3683 VSS.n3682 40.8246
R6597 VSS.n3679 VSS.n3678 40.8246
R6598 VSS.n3675 VSS.n3480 40.8246
R6599 VSS.n3526 VSS.n3519 40.8246
R6600 VSS.n3554 VSS.n3553 40.8246
R6601 VSS.n3550 VSS.n3535 40.8246
R6602 VSS.n3542 VSS.n3541 40.8246
R6603 VSS.n4504 VSS.n1446 40.8246
R6604 VSS.n4573 VSS.n1447 40.8246
R6605 VSS.n4562 VSS.n4561 40.8246
R6606 VSS.n4558 VSS.n4534 40.8246
R6607 VSS.n4547 VSS.n26 40.8246
R6608 VSS.n4546 VSS.n4545 40.8246
R6609 VSS.n4560 VSS.n4559 40.8246
R6610 VSS.n4532 VSS.n4531 40.8246
R6611 VSS.n4575 VSS.n4574 40.8246
R6612 VSS.n4503 VSS.n73 40.8246
R6613 VSS.n3544 VSS.n3543 40.8246
R6614 VSS.n3552 VSS.n3551 40.8246
R6615 VSS.n3534 VSS.n3533 40.8246
R6616 VSS.n3525 VSS.n3524 40.8246
R6617 VSS.n3677 VSS.n3676 40.8246
R6618 VSS.n3475 VSS.n3474 40.8246
R6619 VSS.n3466 VSS.n3465 40.8246
R6620 VSS.n3457 VSS.n3456 40.8246
R6621 VSS.n4880 VSS.n4879 40.8246
R6622 VSS.n970 VSS.n969 40.8246
R6623 VSS.n871 VSS.n848 40.8246
R6624 VSS.n854 VSS.n850 40.8246
R6625 VSS.n853 VSS.n852 40.8246
R6626 VSS.n5133 VSS.n5132 40.8246
R6627 VSS.n432 VSS.n431 40.8246
R6628 VSS.n583 VSS.n569 40.8246
R6629 VSS.n574 VSS.n572 40.8246
R6630 VSS.n5341 VSS.n5340 40.8246
R6631 VSS.n2280 VSS.n177 40.8246
R6632 VSS.n2284 VSS.n2283 40.8246
R6633 VSS.n5429 VSS.n86 40.8246
R6634 VSS.n139 VSS.n88 40.8246
R6635 VSS.n139 VSS.n135 40.8246
R6636 VSS.n143 VSS.n89 40.8246
R6637 VSS.n143 VSS.n136 40.8246
R6638 VSS.n147 VSS.n90 40.8246
R6639 VSS.n147 VSS.n137 40.8246
R6640 VSS.n138 VSS.n91 40.8246
R6641 VSS.n156 VSS.n138 40.8246
R6642 VSS.n152 VSS.n92 40.8246
R6643 VSS.n5427 VSS.n93 40.8246
R6644 VSS.n5425 VSS.n94 40.8246
R6645 VSS.n152 VSS.n93 40.8246
R6646 VSS.n156 VSS.n155 40.8246
R6647 VSS.n155 VSS.n92 40.8246
R6648 VSS.n149 VSS.n137 40.8246
R6649 VSS.n149 VSS.n91 40.8246
R6650 VSS.n145 VSS.n136 40.8246
R6651 VSS.n145 VSS.n90 40.8246
R6652 VSS.n141 VSS.n135 40.8246
R6653 VSS.n141 VSS.n89 40.8246
R6654 VSS.n5432 VSS.n84 40.8246
R6655 VSS.n592 VSS.n80 40.8246
R6656 VSS.n87 VSS.n86 40.8246
R6657 VSS.n88 VSS.n87 40.8246
R6658 VSS.n643 VSS.n642 40.8246
R6659 VSS.n635 VSS.n322 40.8246
R6660 VSS.n5240 VSS.n5239 40.8246
R6661 VSS.n318 VSS.n304 40.8246
R6662 VSS.n316 VSS.n311 40.8246
R6663 VSS.n314 VSS.n305 40.8246
R6664 VSS.n312 VSS.n310 40.8246
R6665 VSS.n5242 VSS.n306 40.8246
R6666 VSS.n5244 VSS.n5243 40.8246
R6667 VSS.n5246 VSS.n307 40.8246
R6668 VSS.n5249 VSS.n308 40.8246
R6669 VSS.n4996 VSS.n4995 40.8246
R6670 VSS.n758 VSS.n744 40.8246
R6671 VSS.n756 VSS.n751 40.8246
R6672 VSS.n754 VSS.n745 40.8246
R6673 VSS.n752 VSS.n750 40.8246
R6674 VSS.n4998 VSS.n746 40.8246
R6675 VSS.n5000 VSS.n4999 40.8246
R6676 VSS.n5002 VSS.n747 40.8246
R6677 VSS.n5005 VSS.n748 40.8246
R6678 VSS.n4407 VSS.n4406 40.8246
R6679 VSS.n1582 VSS.n1568 40.8246
R6680 VSS.n1580 VSS.n1575 40.8246
R6681 VSS.n1578 VSS.n1569 40.8246
R6682 VSS.n1576 VSS.n1574 40.8246
R6683 VSS.n4409 VSS.n1570 40.8246
R6684 VSS.n4411 VSS.n4410 40.8246
R6685 VSS.n4413 VSS.n1571 40.8246
R6686 VSS.n4416 VSS.n1572 40.8246
R6687 VSS.n1256 VSS.n1226 40.8246
R6688 VSS.n1255 VSS.n1254 40.8246
R6689 VSS.n1253 VSS.n1252 40.8246
R6690 VSS.n1251 VSS.n1250 40.8246
R6691 VSS.n1247 VSS.n1230 40.8246
R6692 VSS.n1246 VSS.n1245 40.8246
R6693 VSS.n1244 VSS.n1243 40.8246
R6694 VSS.n1242 VSS.n1241 40.8246
R6695 VSS.n1238 VSS.n1233 40.8246
R6696 VSS.n1237 VSS.n1236 40.8246
R6697 VSS.n1236 VSS.n1235 40.8246
R6698 VSS.n1208 VSS.n1204 40.8246
R6699 VSS.n1238 VSS.n1237 40.8246
R6700 VSS.n1241 VSS.n1233 40.8246
R6701 VSS.n1243 VSS.n1242 40.8246
R6702 VSS.n1245 VSS.n1244 40.8246
R6703 VSS.n1247 VSS.n1246 40.8246
R6704 VSS.n1250 VSS.n1230 40.8246
R6705 VSS.n1252 VSS.n1251 40.8246
R6706 VSS.n1254 VSS.n1253 40.8246
R6707 VSS.n1256 VSS.n1255 40.8246
R6708 VSS.n1226 VSS.n1220 40.8246
R6709 VSS.n4718 VSS.n4717 40.8246
R6710 VSS.n1280 VSS.n1187 40.8246
R6711 VSS.n1281 VSS.n1280 40.8246
R6712 VSS.n1285 VSS.n1188 40.8246
R6713 VSS.n1286 VSS.n1285 40.8246
R6714 VSS.n1290 VSS.n1189 40.8246
R6715 VSS.n1291 VSS.n1290 40.8246
R6716 VSS.n1295 VSS.n1190 40.8246
R6717 VSS.n1296 VSS.n1295 40.8246
R6718 VSS.n1300 VSS.n1191 40.8246
R6719 VSS.n1299 VSS.n1192 40.8246
R6720 VSS.n1300 VSS.n1299 40.8246
R6721 VSS.n1297 VSS.n1296 40.8246
R6722 VSS.n1297 VSS.n1191 40.8246
R6723 VSS.n1292 VSS.n1291 40.8246
R6724 VSS.n1292 VSS.n1190 40.8246
R6725 VSS.n1287 VSS.n1286 40.8246
R6726 VSS.n1287 VSS.n1189 40.8246
R6727 VSS.n1282 VSS.n1281 40.8246
R6728 VSS.n1282 VSS.n1188 40.8246
R6729 VSS.n1337 VSS.n1336 40.8246
R6730 VSS.n1335 VSS.n1334 40.8246
R6731 VSS.n1333 VSS.n1332 40.8246
R6732 VSS.n1329 VSS.n1309 40.8246
R6733 VSS.n1328 VSS.n1327 40.8246
R6734 VSS.n1326 VSS.n1325 40.8246
R6735 VSS.n1324 VSS.n1323 40.8246
R6736 VSS.n1320 VSS.n1312 40.8246
R6737 VSS.n1319 VSS.n1318 40.8246
R6738 VSS.n1317 VSS.n1316 40.8246
R6739 VSS.n1316 VSS.n1315 40.8246
R6740 VSS.n1318 VSS.n1317 40.8246
R6741 VSS.n1320 VSS.n1319 40.8246
R6742 VSS.n1323 VSS.n1312 40.8246
R6743 VSS.n1325 VSS.n1324 40.8246
R6744 VSS.n1327 VSS.n1326 40.8246
R6745 VSS.n1329 VSS.n1328 40.8246
R6746 VSS.n1332 VSS.n1309 40.8246
R6747 VSS.n1334 VSS.n1333 40.8246
R6748 VSS.n1336 VSS.n1335 40.8246
R6749 VSS.n1338 VSS.n1337 40.8246
R6750 VSS.n729 VSS.n725 40.8246
R6751 VSS.n5043 VSS.n5042 40.8246
R6752 VSS.n5039 VSS.n5019 40.8246
R6753 VSS.n5037 VSS.n5018 40.8246
R6754 VSS.n5036 VSS.n5035 40.8246
R6755 VSS.n5023 VSS.n5017 40.8246
R6756 VSS.n5025 VSS.n5021 40.8246
R6757 VSS.n5027 VSS.n5016 40.8246
R6758 VSS.n5029 VSS.n5022 40.8246
R6759 VSS.n5032 VSS.n5015 40.8246
R6760 VSS.n5033 VSS.n5014 40.8246
R6761 VSS.n5033 VSS.n5032 40.8246
R6762 VSS.n5029 VSS.n5015 40.8246
R6763 VSS.n5027 VSS.n5022 40.8246
R6764 VSS.n5025 VSS.n5016 40.8246
R6765 VSS.n5023 VSS.n5021 40.8246
R6766 VSS.n5035 VSS.n5017 40.8246
R6767 VSS.n5037 VSS.n5036 40.8246
R6768 VSS.n5039 VSS.n5018 40.8246
R6769 VSS.n5042 VSS.n5019 40.8246
R6770 VSS.n5286 VSS.n5285 40.8246
R6771 VSS.n5284 VSS.n5283 40.8246
R6772 VSS.n5282 VSS.n5281 40.8246
R6773 VSS.n276 VSS.n271 40.8246
R6774 VSS.n278 VSS.n277 40.8246
R6775 VSS.n5270 VSS.n279 40.8246
R6776 VSS.n5269 VSS.n5268 40.8246
R6777 VSS.n292 VSS.n280 40.8246
R6778 VSS.n294 VSS.n293 40.8246
R6779 VSS.n5257 VSS.n295 40.8246
R6780 VSS.n5256 VSS.n5255 40.8246
R6781 VSS.n5079 VSS.n5078 40.8246
R6782 VSS.n5077 VSS.n5076 40.8246
R6783 VSS.n5075 VSS.n5074 40.8246
R6784 VSS.n704 VSS.n699 40.8246
R6785 VSS.n706 VSS.n705 40.8246
R6786 VSS.n5063 VSS.n707 40.8246
R6787 VSS.n5062 VSS.n5061 40.8246
R6788 VSS.n720 VSS.n708 40.8246
R6789 VSS.n722 VSS.n721 40.8246
R6790 VSS.n5050 VSS.n723 40.8246
R6791 VSS.n5049 VSS.n5048 40.8246
R6792 VSS.n3761 VSS.n3760 40.8246
R6793 VSS.n3763 VSS.n3762 40.8246
R6794 VSS.n3776 VSS.n3764 40.8246
R6795 VSS.n3775 VSS.n3774 40.8246
R6796 VSS.n3773 VSS.n3772 40.8246
R6797 VSS.n3771 VSS.n3770 40.8246
R6798 VSS.n3769 VSS.n3768 40.8246
R6799 VSS.n3767 VSS.n3766 40.8246
R6800 VSS.n3806 VSS.n3755 40.8246
R6801 VSS.n3809 VSS.n3807 40.8246
R6802 VSS.n3808 VSS.n735 40.8246
R6803 VSS.n4453 VSS.n4452 40.8246
R6804 VSS.n4451 VSS.n4450 40.8246
R6805 VSS.n4449 VSS.n4448 40.8246
R6806 VSS.n1541 VSS.n1536 40.8246
R6807 VSS.n1543 VSS.n1542 40.8246
R6808 VSS.n4437 VSS.n1544 40.8246
R6809 VSS.n4436 VSS.n4435 40.8246
R6810 VSS.n1557 VSS.n1545 40.8246
R6811 VSS.n1559 VSS.n1558 40.8246
R6812 VSS.n4424 VSS.n1560 40.8246
R6813 VSS.n4423 VSS.n4422 40.8246
R6814 VSS.n4318 VSS.n4317 40.8246
R6815 VSS.n4316 VSS.n4315 40.8246
R6816 VSS.n4353 VSS.n1758 40.8246
R6817 VSS.n4352 VSS.n4351 40.8246
R6818 VSS.n4350 VSS.n4349 40.8246
R6819 VSS.n2420 VSS.n1760 40.8246
R6820 VSS.n2419 VSS.n2418 40.8246
R6821 VSS.n2417 VSS.n2416 40.8246
R6822 VSS.n2415 VSS.n2414 40.8246
R6823 VSS.n2512 VSS.n2410 40.8246
R6824 VSS.n2514 VSS.n2513 40.8246
R6825 VSS.n4027 VSS.n4012 40.8246
R6826 VSS.n4026 VSS.n4016 40.8246
R6827 VSS.n4038 VSS.n4037 40.8246
R6828 VSS.n4034 VSS.n4017 40.8246
R6829 VSS.n4032 VSS.n4025 40.8246
R6830 VSS.n4030 VSS.n4018 40.8246
R6831 VSS.n4024 VSS.n4023 40.8246
R6832 VSS.n4041 VSS.n4019 40.8246
R6833 VSS.n4040 VSS.n4020 40.8246
R6834 VSS.n4046 VSS.n4045 40.8246
R6835 VSS.n4045 VSS.n4021 40.8246
R6836 VSS.n4046 VSS.n4020 40.8246
R6837 VSS.n4041 VSS.n4040 40.8246
R6838 VSS.n4023 VSS.n4019 40.8246
R6839 VSS.n4030 VSS.n4024 40.8246
R6840 VSS.n4032 VSS.n4018 40.8246
R6841 VSS.n4034 VSS.n4025 40.8246
R6842 VSS.n4037 VSS.n4017 40.8246
R6843 VSS.n4038 VSS.n4026 40.8246
R6844 VSS.n4027 VSS.n4016 40.8246
R6845 VSS.n4048 VSS.n4012 40.8246
R6846 VSS.n1163 VSS.n1159 40.8246
R6847 VSS.n3902 VSS.n3901 40.8246
R6848 VSS.n3898 VSS.n3872 40.8246
R6849 VSS.n3897 VSS.n3896 40.8246
R6850 VSS.n3895 VSS.n3894 40.8246
R6851 VSS.n3893 VSS.n3892 40.8246
R6852 VSS.n3889 VSS.n3875 40.8246
R6853 VSS.n3888 VSS.n3887 40.8246
R6854 VSS.n3886 VSS.n3885 40.8246
R6855 VSS.n3884 VSS.n3883 40.8246
R6856 VSS.n3880 VSS.n3878 40.8246
R6857 VSS.n3880 VSS.n3879 40.8246
R6858 VSS.n3883 VSS.n3878 40.8246
R6859 VSS.n3885 VSS.n3884 40.8246
R6860 VSS.n3887 VSS.n3886 40.8246
R6861 VSS.n3889 VSS.n3888 40.8246
R6862 VSS.n3892 VSS.n3875 40.8246
R6863 VSS.n3894 VSS.n3893 40.8246
R6864 VSS.n3896 VSS.n3895 40.8246
R6865 VSS.n3898 VSS.n3897 40.8246
R6866 VSS.n3901 VSS.n3872 40.8246
R6867 VSS.n3903 VSS.n3902 40.8246
R6868 VSS.n2713 VSS.n1266 40.8246
R6869 VSS.n2715 VSS.n2714 40.8246
R6870 VSS.n2082 VSS.n1267 40.8246
R6871 VSS.n2084 VSS.n2083 40.8246
R6872 VSS.n2228 VSS.n1268 40.8246
R6873 VSS.n2227 VSS.n2226 40.8246
R6874 VSS.n2093 VSS.n1269 40.8246
R6875 VSS.n2095 VSS.n2094 40.8246
R6876 VSS.n2211 VSS.n1270 40.8246
R6877 VSS.n2210 VSS.n1259 40.8246
R6878 VSS.n4685 VSS.n4684 40.8246
R6879 VSS.n3019 VSS.n1222 40.8246
R6880 VSS.n3021 VSS.n3020 40.8246
R6881 VSS.n2859 VSS.n1271 40.8246
R6882 VSS.n2861 VSS.n2860 40.8246
R6883 VSS.n3006 VSS.n1272 40.8246
R6884 VSS.n3005 VSS.n3004 40.8246
R6885 VSS.n2870 VSS.n1273 40.8246
R6886 VSS.n2872 VSS.n2871 40.8246
R6887 VSS.n2989 VSS.n1274 40.8246
R6888 VSS.n2988 VSS.n2987 40.8246
R6889 VSS.n1342 VSS.n1341 40.8246
R6890 VSS.n4790 VSS.n1059 40.8246
R6891 VSS.n4789 VSS.n4788 40.8246
R6892 VSS.n1343 VSS.n1061 40.8246
R6893 VSS.n1345 VSS.n1344 40.8246
R6894 VSS.n3844 VSS.n1346 40.8246
R6895 VSS.n3846 VSS.n3845 40.8246
R6896 VSS.n3853 VSS.n1347 40.8246
R6897 VSS.n3855 VSS.n3854 40.8246
R6898 VSS.n3862 VSS.n1348 40.8246
R6899 VSS.n3864 VSS.n3863 40.8246
R6900 VSS.n3922 VSS.n1349 40.8246
R6901 VSS.n3927 VSS.n1350 40.8246
R6902 VSS.n3929 VSS.n3928 40.8246
R6903 VSS.n3282 VSS.n1351 40.8246
R6904 VSS.n3284 VSS.n3283 40.8246
R6905 VSS.n3403 VSS.n1352 40.8246
R6906 VSS.n3402 VSS.n3401 40.8246
R6907 VSS.n3293 VSS.n1353 40.8246
R6908 VSS.n3295 VSS.n3294 40.8246
R6909 VSS.n3386 VSS.n1354 40.8246
R6910 VSS.n3385 VSS.n3384 40.8246
R6911 VSS.n4011 VSS.n1355 40.8246
R6912 VSS.n4294 VSS.n1264 40.8246
R6913 VSS.n4293 VSS.n4292 40.8246
R6914 VSS.n1786 VSS.n1263 40.8246
R6915 VSS.n1788 VSS.n1787 40.8246
R6916 VSS.n2466 VSS.n1262 40.8246
R6917 VSS.n2468 VSS.n2467 40.8246
R6918 VSS.n2475 VSS.n1261 40.8246
R6919 VSS.n2477 VSS.n2476 40.8246
R6920 VSS.n2483 VSS.n1260 40.8246
R6921 VSS.n2482 VSS.n1356 40.8246
R6922 VSS.n4682 VSS.n4681 40.8246
R6923 VSS.n2708 VSS.n1266 40.8246
R6924 VSS.n2715 VSS.n1267 40.8246
R6925 VSS.n2084 VSS.n1268 40.8246
R6926 VSS.n2226 VSS.n1269 40.8246
R6927 VSS.n2095 VSS.n1270 40.8246
R6928 VSS.n4684 VSS.n1259 40.8246
R6929 VSS.n4687 VSS.n1222 40.8246
R6930 VSS.n3021 VSS.n1271 40.8246
R6931 VSS.n2861 VSS.n1272 40.8246
R6932 VSS.n3004 VSS.n1273 40.8246
R6933 VSS.n2872 VSS.n1274 40.8246
R6934 VSS.n2987 VSS.n1342 40.8246
R6935 VSS.n1277 VSS.n1059 40.8246
R6936 VSS.n4788 VSS.n1061 40.8246
R6937 VSS.n1346 VSS.n1345 40.8246
R6938 VSS.n3846 VSS.n1347 40.8246
R6939 VSS.n3855 VSS.n1348 40.8246
R6940 VSS.n3864 VSS.n1349 40.8246
R6941 VSS.n3868 VSS.n1350 40.8246
R6942 VSS.n3929 VSS.n1351 40.8246
R6943 VSS.n3284 VSS.n1352 40.8246
R6944 VSS.n3401 VSS.n1353 40.8246
R6945 VSS.n3295 VSS.n1354 40.8246
R6946 VSS.n3384 VSS.n1355 40.8246
R6947 VSS.n4013 VSS.n1264 40.8246
R6948 VSS.n3386 VSS.n3385 40.8246
R6949 VSS.n3294 VSS.n3293 40.8246
R6950 VSS.n3403 VSS.n3402 40.8246
R6951 VSS.n3283 VSS.n3282 40.8246
R6952 VSS.n3928 VSS.n3927 40.8246
R6953 VSS.n3863 VSS.n3862 40.8246
R6954 VSS.n3854 VSS.n3853 40.8246
R6955 VSS.n3845 VSS.n3844 40.8246
R6956 VSS.n1344 VSS.n1343 40.8246
R6957 VSS.n4790 VSS.n4789 40.8246
R6958 VSS.n2989 VSS.n2988 40.8246
R6959 VSS.n2871 VSS.n2870 40.8246
R6960 VSS.n3006 VSS.n3005 40.8246
R6961 VSS.n2860 VSS.n2859 40.8246
R6962 VSS.n3020 VSS.n3019 40.8246
R6963 VSS.n2211 VSS.n2210 40.8246
R6964 VSS.n2094 VSS.n2093 40.8246
R6965 VSS.n2228 VSS.n2227 40.8246
R6966 VSS.n2083 VSS.n2082 40.8246
R6967 VSS.n2714 VSS.n2713 40.8246
R6968 VSS.n3097 VSS.n3066 40.8246
R6969 VSS.n3076 VSS.n3067 40.8246
R6970 VSS.n3076 VSS.n3074 40.8246
R6971 VSS.n3080 VSS.n3068 40.8246
R6972 VSS.n3080 VSS.n3075 40.8246
R6973 VSS.n3085 VSS.n3069 40.8246
R6974 VSS.n3087 VSS.n3085 40.8246
R6975 VSS.n3090 VSS.n3070 40.8246
R6976 VSS.n3090 VSS.n3089 40.8246
R6977 VSS.n3095 VSS.n3094 40.8246
R6978 VSS.n3072 VSS.n1195 40.8246
R6979 VSS.n3094 VSS.n3072 40.8246
R6980 VSS.n3089 VSS.n3071 40.8246
R6981 VSS.n3095 VSS.n3071 40.8246
R6982 VSS.n3087 VSS.n3086 40.8246
R6983 VSS.n3086 VSS.n3070 40.8246
R6984 VSS.n3082 VSS.n3075 40.8246
R6985 VSS.n3082 VSS.n3069 40.8246
R6986 VSS.n3078 VSS.n3074 40.8246
R6987 VSS.n3078 VSS.n3068 40.8246
R6988 VSS.n3182 VSS.n3152 40.8246
R6989 VSS.n3161 VSS.n3153 40.8246
R6990 VSS.n3161 VSS.n3158 40.8246
R6991 VSS.n3165 VSS.n3154 40.8246
R6992 VSS.n3165 VSS.n3159 40.8246
R6993 VSS.n3169 VSS.n3155 40.8246
R6994 VSS.n3169 VSS.n3160 40.8246
R6995 VSS.n3175 VSS.n3156 40.8246
R6996 VSS.n3176 VSS.n3175 40.8246
R6997 VSS.n3180 VSS.n3179 40.8246
R6998 VSS.n3178 VSS.n1160 40.8246
R6999 VSS.n3179 VSS.n3178 40.8246
R7000 VSS.n3176 VSS.n3157 40.8246
R7001 VSS.n3180 VSS.n3157 40.8246
R7002 VSS.n3171 VSS.n3160 40.8246
R7003 VSS.n3171 VSS.n3156 40.8246
R7004 VSS.n3167 VSS.n3159 40.8246
R7005 VSS.n3167 VSS.n3155 40.8246
R7006 VSS.n3163 VSS.n3158 40.8246
R7007 VSS.n3163 VSS.n3154 40.8246
R7008 VSS.n4076 VSS.n1914 40.8246
R7009 VSS.n3980 VSS.n1916 40.8246
R7010 VSS.n3980 VSS.n3976 40.8246
R7011 VSS.n3984 VSS.n1917 40.8246
R7012 VSS.n3984 VSS.n3977 40.8246
R7013 VSS.n3978 VSS.n1918 40.8246
R7014 VSS.n3991 VSS.n3978 40.8246
R7015 VSS.n3975 VSS.n1919 40.8246
R7016 VSS.n3993 VSS.n3975 40.8246
R7017 VSS.n3996 VSS.n1920 40.8246
R7018 VSS.n4074 VSS.n1921 40.8246
R7019 VSS.n3996 VSS.n1921 40.8246
R7020 VSS.n3994 VSS.n3993 40.8246
R7021 VSS.n3994 VSS.n1920 40.8246
R7022 VSS.n3991 VSS.n3990 40.8246
R7023 VSS.n3990 VSS.n1919 40.8246
R7024 VSS.n3986 VSS.n3977 40.8246
R7025 VSS.n3986 VSS.n1918 40.8246
R7026 VSS.n3982 VSS.n3976 40.8246
R7027 VSS.n3982 VSS.n1917 40.8246
R7028 VSS.n4000 VSS.n3999 40.8246
R7029 VSS.n2680 VSS.n2679 40.8246
R7030 VSS.n2745 VSS.n2066 40.8246
R7031 VSS.n2744 VSS.n2743 40.8246
R7032 VSS.n2133 VSS.n2067 40.8246
R7033 VSS.n2132 VSS.n2131 40.8246
R7034 VSS.n2130 VSS.n2129 40.8246
R7035 VSS.n2152 VSS.n2126 40.8246
R7036 VSS.n2154 VSS.n2153 40.8246
R7037 VSS.n2156 VSS.n2155 40.8246
R7038 VSS.n2159 VSS.n2157 40.8246
R7039 VSS.n2158 VSS.n1201 40.8246
R7040 VSS.n2846 VSS.n2845 40.8246
R7041 VSS.n3051 VSS.n2023 40.8246
R7042 VSS.n3050 VSS.n3049 40.8246
R7043 VSS.n2912 VSS.n2024 40.8246
R7044 VSS.n2911 VSS.n2910 40.8246
R7045 VSS.n2909 VSS.n2908 40.8246
R7046 VSS.n2931 VSS.n2905 40.8246
R7047 VSS.n2933 VSS.n2932 40.8246
R7048 VSS.n2935 VSS.n2934 40.8246
R7049 VSS.n2938 VSS.n2936 40.8246
R7050 VSS.n2937 VSS.n1197 40.8246
R7051 VSS.n4765 VSS.n4764 40.8246
R7052 VSS.n4763 VSS.n4762 40.8246
R7053 VSS.n4761 VSS.n4760 40.8246
R7054 VSS.n1138 VSS.n1133 40.8246
R7055 VSS.n1140 VSS.n1139 40.8246
R7056 VSS.n4749 VSS.n1141 40.8246
R7057 VSS.n4748 VSS.n4747 40.8246
R7058 VSS.n1154 VSS.n1142 40.8246
R7059 VSS.n1156 VSS.n1155 40.8246
R7060 VSS.n4736 VSS.n1157 40.8246
R7061 VSS.n4735 VSS.n4734 40.8246
R7062 VSS.n3269 VSS.n3268 40.8246
R7063 VSS.n3959 VSS.n1947 40.8246
R7064 VSS.n3958 VSS.n3957 40.8246
R7065 VSS.n3315 VSS.n1948 40.8246
R7066 VSS.n3314 VSS.n3313 40.8246
R7067 VSS.n3312 VSS.n3311 40.8246
R7068 VSS.n3334 VSS.n3308 40.8246
R7069 VSS.n3336 VSS.n3335 40.8246
R7070 VSS.n3338 VSS.n3337 40.8246
R7071 VSS.n3968 VSS.n1923 40.8246
R7072 VSS.n3970 VSS.n3969 40.8246
R7073 VSS.n4255 VSS.n1837 40.8246
R7074 VSS.n4254 VSS.n4253 40.8246
R7075 VSS.n4252 VSS.n4251 40.8246
R7076 VSS.n4250 VSS.n4249 40.8246
R7077 VSS.n4248 VSS.n4247 40.8246
R7078 VSS.n4237 VSS.n1841 40.8246
R7079 VSS.n4236 VSS.n4235 40.8246
R7080 VSS.n4225 VSS.n1843 40.8246
R7081 VSS.n4224 VSS.n4223 40.8246
R7082 VSS.n4216 VSS.n1847 40.8246
R7083 VSS.n4215 VSS.n4214 40.8246
R7084 VSS.n2760 VSS.n2037 40.8246
R7085 VSS.n2790 VSS.n2760 40.8246
R7086 VSS.n3066 VSS.n1994 40.8246
R7087 VSS.n3067 VSS.n1994 40.8246
R7088 VSS.n3152 VSS.n1960 40.8246
R7089 VSS.n3153 VSS.n1960 40.8246
R7090 VSS.n1915 VSS.n1914 40.8246
R7091 VSS.n1916 VSS.n1915 40.8246
R7092 VSS.n2679 VSS.n2066 40.8246
R7093 VSS.n2743 VSS.n2067 40.8246
R7094 VSS.n2131 VSS.n2130 40.8246
R7095 VSS.n2153 VSS.n2152 40.8246
R7096 VSS.n2157 VSS.n2156 40.8246
R7097 VSS.n2846 VSS.n2023 40.8246
R7098 VSS.n3049 VSS.n2024 40.8246
R7099 VSS.n2910 VSS.n2909 40.8246
R7100 VSS.n2932 VSS.n2931 40.8246
R7101 VSS.n2936 VSS.n2935 40.8246
R7102 VSS.n4764 VSS.n4763 40.8246
R7103 VSS.n4760 VSS.n1133 40.8246
R7104 VSS.n1141 VSS.n1140 40.8246
R7105 VSS.n4747 VSS.n1142 40.8246
R7106 VSS.n1157 VSS.n1156 40.8246
R7107 VSS.n3269 VSS.n1947 40.8246
R7108 VSS.n3957 VSS.n1948 40.8246
R7109 VSS.n3313 VSS.n3312 40.8246
R7110 VSS.n3335 VSS.n3334 40.8246
R7111 VSS.n3338 VSS.n1923 40.8246
R7112 VSS.n4255 VSS.n4254 40.8246
R7113 VSS.n4251 VSS.n4250 40.8246
R7114 VSS.n4247 VSS.n1841 40.8246
R7115 VSS.n4235 VSS.n1843 40.8246
R7116 VSS.n4223 VSS.n1847 40.8246
R7117 VSS.n4216 VSS.n4215 40.8246
R7118 VSS.n4225 VSS.n4224 40.8246
R7119 VSS.n4237 VSS.n4236 40.8246
R7120 VSS.n4249 VSS.n4248 40.8246
R7121 VSS.n4253 VSS.n4252 40.8246
R7122 VSS.n1837 VSS.n1836 40.8246
R7123 VSS.n3969 VSS.n3968 40.8246
R7124 VSS.n3337 VSS.n3336 40.8246
R7125 VSS.n3311 VSS.n3308 40.8246
R7126 VSS.n3315 VSS.n3314 40.8246
R7127 VSS.n3959 VSS.n3958 40.8246
R7128 VSS.n3268 VSS.n3267 40.8246
R7129 VSS.n4736 VSS.n4735 40.8246
R7130 VSS.n1155 VSS.n1154 40.8246
R7131 VSS.n4749 VSS.n4748 40.8246
R7132 VSS.n1139 VSS.n1138 40.8246
R7133 VSS.n4762 VSS.n4761 40.8246
R7134 VSS.n4766 VSS.n4765 40.8246
R7135 VSS.n2938 VSS.n2937 40.8246
R7136 VSS.n2934 VSS.n2933 40.8246
R7137 VSS.n2908 VSS.n2905 40.8246
R7138 VSS.n2912 VSS.n2911 40.8246
R7139 VSS.n3051 VSS.n3050 40.8246
R7140 VSS.n2845 VSS.n2844 40.8246
R7141 VSS.n2159 VSS.n2158 40.8246
R7142 VSS.n2155 VSS.n2154 40.8246
R7143 VSS.n2129 VSS.n2126 40.8246
R7144 VSS.n2133 VSS.n2132 40.8246
R7145 VSS.n2745 VSS.n2744 40.8246
R7146 VSS.n2681 VSS.n2680 40.8246
R7147 VSS.n4708 VSS.n1204 40.8246
R7148 VSS.n4717 VSS.n4716 40.8246
R7149 VSS.n4716 VSS.n1187 40.8246
R7150 VSS.n4729 VSS.n1159 40.8246
R7151 VSS.n4072 VSS.n4000 40.8246
R7152 VSS.n4292 VSS.n1263 40.8246
R7153 VSS.n1788 VSS.n1262 40.8246
R7154 VSS.n2468 VSS.n1261 40.8246
R7155 VSS.n2477 VSS.n1260 40.8246
R7156 VSS.n4682 VSS.n1356 40.8246
R7157 VSS.n2483 VSS.n2482 40.8246
R7158 VSS.n2476 VSS.n2475 40.8246
R7159 VSS.n2467 VSS.n2466 40.8246
R7160 VSS.n1787 VSS.n1786 40.8246
R7161 VSS.n4294 VSS.n4293 40.8246
R7162 VSS.n1235 VSS.n298 40.8246
R7163 VSS.n1315 VSS.n726 40.8246
R7164 VSS.n3879 VSS.n739 40.8246
R7165 VSS.n4021 VSS.n1562 40.8246
R7166 VSS.n5285 VSS.n5284 40.8246
R7167 VSS.n5281 VSS.n271 40.8246
R7168 VSS.n279 VSS.n278 40.8246
R7169 VSS.n5268 VSS.n280 40.8246
R7170 VSS.n295 VSS.n294 40.8246
R7171 VSS.n5078 VSS.n5077 40.8246
R7172 VSS.n5074 VSS.n699 40.8246
R7173 VSS.n707 VSS.n706 40.8246
R7174 VSS.n5061 VSS.n708 40.8246
R7175 VSS.n723 VSS.n722 40.8246
R7176 VSS.n3762 VSS.n3761 40.8246
R7177 VSS.n3776 VSS.n3775 40.8246
R7178 VSS.n3772 VSS.n3771 40.8246
R7179 VSS.n3768 VSS.n3767 40.8246
R7180 VSS.n3807 VSS.n3806 40.8246
R7181 VSS.n4452 VSS.n4451 40.8246
R7182 VSS.n4448 VSS.n1536 40.8246
R7183 VSS.n1544 VSS.n1543 40.8246
R7184 VSS.n4435 VSS.n1545 40.8246
R7185 VSS.n1560 VSS.n1559 40.8246
R7186 VSS.n4317 VSS.n4316 40.8246
R7187 VSS.n4353 VSS.n4352 40.8246
R7188 VSS.n4349 VSS.n1760 40.8246
R7189 VSS.n2418 VSS.n2417 40.8246
R7190 VSS.n2414 VSS.n2410 40.8246
R7191 VSS.n2513 VSS.n2512 40.8246
R7192 VSS.n2416 VSS.n2415 40.8246
R7193 VSS.n2420 VSS.n2419 40.8246
R7194 VSS.n4351 VSS.n4350 40.8246
R7195 VSS.n4315 VSS.n1758 40.8246
R7196 VSS.n4319 VSS.n4318 40.8246
R7197 VSS.n4424 VSS.n4423 40.8246
R7198 VSS.n1558 VSS.n1557 40.8246
R7199 VSS.n4437 VSS.n4436 40.8246
R7200 VSS.n1542 VSS.n1541 40.8246
R7201 VSS.n4450 VSS.n4449 40.8246
R7202 VSS.n4454 VSS.n4453 40.8246
R7203 VSS.n3809 VSS.n3808 40.8246
R7204 VSS.n3766 VSS.n3755 40.8246
R7205 VSS.n3770 VSS.n3769 40.8246
R7206 VSS.n3774 VSS.n3773 40.8246
R7207 VSS.n3764 VSS.n3763 40.8246
R7208 VSS.n3760 VSS.n731 40.8246
R7209 VSS.n5050 VSS.n5049 40.8246
R7210 VSS.n721 VSS.n720 40.8246
R7211 VSS.n5063 VSS.n5062 40.8246
R7212 VSS.n705 VSS.n704 40.8246
R7213 VSS.n5076 VSS.n5075 40.8246
R7214 VSS.n5080 VSS.n5079 40.8246
R7215 VSS.n5257 VSS.n5256 40.8246
R7216 VSS.n293 VSS.n292 40.8246
R7217 VSS.n5270 VSS.n5269 40.8246
R7218 VSS.n277 VSS.n276 40.8246
R7219 VSS.n5283 VSS.n5282 40.8246
R7220 VSS.n5287 VSS.n5286 40.8246
R7221 VSS.n5250 VSS.n297 40.8246
R7222 VSS.n5252 VSS.n301 40.8246
R7223 VSS.n5043 VSS.n725 40.8246
R7224 VSS.n5045 VSS.n729 40.8246
R7225 VSS.n5006 VSS.n738 40.8246
R7226 VSS.n5008 VSS.n741 40.8246
R7227 VSS.n4417 VSS.n1561 40.8246
R7228 VSS.n4419 VSS.n1565 40.8246
R7229 VSS.n1731 VSS.n1389 40.8246
R7230 VSS.n5535 VSS.n5534 40.8246
R7231 VSS.n5427 VSS.n94 40.8246
R7232 VSS.n5214 VSS.n368 40.8246
R7233 VSS.n4961 VSS.n783 40.8246
R7234 VSS.n5463 VSS.n59 40.8246
R7235 VSS.n5465 VSS.n5464 40.8246
R7236 VSS.n5460 VSS.n64 40.8246
R7237 VSS.n5461 VSS.n5459 40.8246
R7238 VSS.n5456 VSS.n69 40.8246
R7239 VSS.n5454 VSS.n68 40.8246
R7240 VSS.n5453 VSS.n5452 40.8246
R7241 VSS.n5449 VSS.n67 40.8246
R7242 VSS.n5448 VSS.n5447 40.8246
R7243 VSS.n5444 VSS.n66 40.8246
R7244 VSS.n5443 VSS.n5442 40.8246
R7245 VSS.n5439 VSS.n65 40.8246
R7246 VSS.n4657 VSS.n4656 38.5594
R7247 VSS.t12 VSS.t28 38.3242
R7248 VSS.n5234 VSS.t40 36.9872
R7249 VSS.n4641 VSS.n209 36.9872
R7250 VSS.n5436 VSS.t44 36.9872
R7251 VSS.n23 VSS.n20 36.9872
R7252 VSS.n5011 VSS.t31 36.9872
R7253 VSS.n2545 VSS.n269 36.9872
R7254 VSS.n4713 VSS.t38 36.9872
R7255 VSS.n4180 VSS.n1131 36.9872
R7256 VSS.t33 VSS.n1182 36.9872
R7257 VSS.n4683 VSS.n1265 36.9872
R7258 VSS.n1374 VSS.n1369 36.563
R7259 VSS.t8 VSS.n1369 36.563
R7260 VSS.n1402 VSS.n1399 36.563
R7261 VSS.n1872 VSS.n1402 36.563
R7262 VSS.n4641 VSS.n211 34.8534
R7263 VSS.n25 VSS.n20 34.8534
R7264 VSS.n2545 VSS.n270 34.8534
R7265 VSS.n4180 VSS.n1132 34.8534
R7266 VSS.n1265 VSS.n1060 34.8534
R7267 VSS.t79 VSS.n4617 34.7088
R7268 VSS.n4659 VSS.n4658 34.4123
R7269 VSS.n4658 VSS.n4657 34.4123
R7270 VSS.n4663 VSS.n4662 34.4123
R7271 VSS.n4664 VSS.n4663 34.4123
R7272 VSS.n4625 VSS.n4624 34.4123
R7273 VSS.t14 VSS.n4625 34.4123
R7274 VSS.n4627 VSS.n4626 34.4123
R7275 VSS.n4626 VSS.t14 34.4123
R7276 VSS.n4639 VSS.n4638 34.4123
R7277 VSS.t6 VSS.n4639 34.4123
R7278 VSS.n1395 VSS.n1393 34.4123
R7279 VSS.n1873 VSS.n1393 34.4123
R7280 VSS.t13 VSS.t2 32.5395
R7281 VSS.n4419 VSS.n1564 31.2084
R7282 VSS.n5252 VSS.n300 31.2084
R7283 VSS.n676 VSS.n323 31.2084
R7284 VSS.n334 VSS.n330 31.2084
R7285 VSS.n5217 VSS.n5216 31.2084
R7286 VSS.n4964 VSS.n4963 31.2084
R7287 VSS.n5008 VSS.n736 31.2084
R7288 VSS.n4987 VSS.n764 31.2084
R7289 VSS.n1685 VSS.n1653 31.2084
R7290 VSS.n5439 VSS.n5438 31.2084
R7291 VSS.n5429 VSS.n81 31.2084
R7292 VSS.n4689 VSS.n1220 31.2084
R7293 VSS.n4708 VSS.n1202 31.2084
R7294 VSS.n4718 VSS.n1193 31.2084
R7295 VSS.n1338 VSS.n1305 31.2084
R7296 VSS.n5045 VSS.n728 31.2084
R7297 VSS.n4049 VSS.n4048 31.2084
R7298 VSS.n4729 VSS.n1166 31.2084
R7299 VSS.n3904 VSS.n3903 31.2084
R7300 VSS.n4072 VSS.n3973 31.2084
R7301 VSS.n4665 VSS.n4664 25.7064
R7302 VSS.t6 VSS.n1392 25.7064
R7303 VSS.n5212 VSS.n397 24.3817
R7304 VSS.n4959 VSS.n812 24.3817
R7305 VSS.n5473 VSS.n58 24.3817
R7306 VSS.n5425 VSS.n98 24.3817
R7307 VSS.t63 VSS.t85 24.1442
R7308 VSS.n4657 VSS.t40 23.5643
R7309 VSS.n0 VSS.t27 21.5736
R7310 VSS.n4632 VSS.t5 21.5736
R7311 VSS.n1396 VSS.t1 21.5546
R7312 VSS.n4635 VSS.t26 21.4809
R7313 VSS.n1396 VSS.t4 21.4809
R7314 VSS.n1889 VSS.n1888 18.261
R7315 VSS.n2357 VSS.n2339 17.4227
R7316 VSS.n5234 VSS.n209 16.36
R7317 VSS.n5436 VSS.n23 16.36
R7318 VSS.n5011 VSS.n269 16.36
R7319 VSS.n4713 VSS.n1131 16.36
R7320 VSS.n4683 VSS.n1182 16.36
R7321 VSS.n2437 VSS.n2436 16.0005
R7322 VSS.n2440 VSS.n2437 16.0005
R7323 VSS.n2441 VSS.n2440 16.0005
R7324 VSS.n2444 VSS.n2441 16.0005
R7325 VSS.n2445 VSS.n2444 16.0005
R7326 VSS.n2448 VSS.n2445 16.0005
R7327 VSS.n2449 VSS.n2448 16.0005
R7328 VSS.n2452 VSS.n2449 16.0005
R7329 VSS.n4147 VSS.n4145 16.0005
R7330 VSS.n4145 VSS.n4142 16.0005
R7331 VSS.n4142 VSS.n4141 16.0005
R7332 VSS.n4141 VSS.n4138 16.0005
R7333 VSS.n4138 VSS.n4137 16.0005
R7334 VSS.n4137 VSS.n4134 16.0005
R7335 VSS.n4134 VSS.n4133 16.0005
R7336 VSS.n4133 VSS.n4130 16.0005
R7337 VSS.n4094 VSS.n4093 16.0005
R7338 VSS.n4093 VSS.n4090 16.0005
R7339 VSS.n4090 VSS.n4089 16.0005
R7340 VSS.n4089 VSS.n4086 16.0005
R7341 VSS.n4086 VSS.n4085 16.0005
R7342 VSS.n4085 VSS.n4082 16.0005
R7343 VSS.n4082 VSS.n1832 16.0005
R7344 VSS.n4274 VSS.n1832 16.0005
R7345 VSS.n3219 VSS.n3217 16.0005
R7346 VSS.n3217 VSS.n3214 16.0005
R7347 VSS.n3214 VSS.n3213 16.0005
R7348 VSS.n3213 VSS.n3210 16.0005
R7349 VSS.n3210 VSS.n3209 16.0005
R7350 VSS.n3209 VSS.n3206 16.0005
R7351 VSS.n3206 VSS.n3205 16.0005
R7352 VSS.n3205 VSS.n3203 16.0005
R7353 VSS.n3252 VSS.n3251 16.0005
R7354 VSS.n3255 VSS.n3252 16.0005
R7355 VSS.n3256 VSS.n3255 16.0005
R7356 VSS.n3259 VSS.n3256 16.0005
R7357 VSS.n3260 VSS.n3259 16.0005
R7358 VSS.n3263 VSS.n3260 16.0005
R7359 VSS.n3265 VSS.n3263 16.0005
R7360 VSS.n3266 VSS.n3265 16.0005
R7361 VSS.n1978 VSS.n1976 16.0005
R7362 VSS.n1976 VSS.n1973 16.0005
R7363 VSS.n1973 VSS.n1972 16.0005
R7364 VSS.n1972 VSS.n1969 16.0005
R7365 VSS.n1969 VSS.n1968 16.0005
R7366 VSS.n1968 VSS.n1965 16.0005
R7367 VSS.n1965 VSS.n1964 16.0005
R7368 VSS.n1964 VSS.n1961 16.0005
R7369 VSS.n3109 VSS.n3106 16.0005
R7370 VSS.n3106 VSS.n3103 16.0005
R7371 VSS.n3103 VSS.n3102 16.0005
R7372 VSS.n3102 VSS.n3099 16.0005
R7373 VSS.n3099 VSS.n1112 16.0005
R7374 VSS.n4772 VSS.n1112 16.0005
R7375 VSS.n4772 VSS.n4771 16.0005
R7376 VSS.n4771 VSS.n4770 16.0005
R7377 VSS.n2884 VSS.n2883 16.0005
R7378 VSS.n2887 VSS.n2884 16.0005
R7379 VSS.n2888 VSS.n2887 16.0005
R7380 VSS.n2891 VSS.n2888 16.0005
R7381 VSS.n2892 VSS.n2891 16.0005
R7382 VSS.n2895 VSS.n2892 16.0005
R7383 VSS.n2896 VSS.n2895 16.0005
R7384 VSS.n2899 VSS.n2896 16.0005
R7385 VSS.n2829 VSS.n2828 16.0005
R7386 VSS.n2832 VSS.n2829 16.0005
R7387 VSS.n2833 VSS.n2832 16.0005
R7388 VSS.n2836 VSS.n2833 16.0005
R7389 VSS.n2837 VSS.n2836 16.0005
R7390 VSS.n2840 VSS.n2837 16.0005
R7391 VSS.n2842 VSS.n2840 16.0005
R7392 VSS.n2843 VSS.n2842 16.0005
R7393 VSS.n4843 VSS.n4793 16.0005
R7394 VSS.n4843 VSS.n4842 16.0005
R7395 VSS.n4842 VSS.n4841 16.0005
R7396 VSS.n4841 VSS.n4838 16.0005
R7397 VSS.n4838 VSS.n4837 16.0005
R7398 VSS.n4837 VSS.n4834 16.0005
R7399 VSS.n4834 VSS.n4833 16.0005
R7400 VSS.n4833 VSS.n4830 16.0005
R7401 VSS.n1128 VSS.n1127 16.0005
R7402 VSS.n1127 VSS.n1124 16.0005
R7403 VSS.n1124 VSS.n1123 16.0005
R7404 VSS.n1123 VSS.n1120 16.0005
R7405 VSS.n1120 VSS.n1119 16.0005
R7406 VSS.n1119 VSS.n1116 16.0005
R7407 VSS.n1116 VSS.n1115 16.0005
R7408 VSS.n1115 VSS.n1055 16.0005
R7409 VSS.n3417 VSS.n3416 16.0005
R7410 VSS.n3420 VSS.n3417 16.0005
R7411 VSS.n3421 VSS.n3420 16.0005
R7412 VSS.n3424 VSS.n3421 16.0005
R7413 VSS.n3425 VSS.n3424 16.0005
R7414 VSS.n3428 VSS.n3425 16.0005
R7415 VSS.n3429 VSS.n3428 16.0005
R7416 VSS.n3432 VSS.n3429 16.0005
R7417 VSS.n3829 VSS.n3827 16.0005
R7418 VSS.n3827 VSS.n3824 16.0005
R7419 VSS.n3824 VSS.n3823 16.0005
R7420 VSS.n3823 VSS.n3820 16.0005
R7421 VSS.n3820 VSS.n3819 16.0005
R7422 VSS.n3819 VSS.n3816 16.0005
R7423 VSS.n3816 VSS.n3815 16.0005
R7424 VSS.n3815 VSS.n3812 16.0005
R7425 VSS.n2340 VSS.n266 16.0005
R7426 VSS.n2343 VSS.n2340 16.0005
R7427 VSS.n2344 VSS.n2343 16.0005
R7428 VSS.n2347 VSS.n2344 16.0005
R7429 VSS.n2348 VSS.n2347 16.0005
R7430 VSS.n2351 VSS.n2348 16.0005
R7431 VSS.n2352 VSS.n2351 16.0005
R7432 VSS.n2355 VSS.n2352 16.0005
R7433 VSS.n535 VSS.n534 16.0005
R7434 VSS.n538 VSS.n535 16.0005
R7435 VSS.n539 VSS.n538 16.0005
R7436 VSS.n542 VSS.n539 16.0005
R7437 VSS.n543 VSS.n542 16.0005
R7438 VSS.n546 VSS.n543 16.0005
R7439 VSS.n547 VSS.n546 16.0005
R7440 VSS.n550 VSS.n547 16.0005
R7441 VSS.n5353 VSS.n5352 16.0005
R7442 VSS.n5356 VSS.n5353 16.0005
R7443 VSS.n5357 VSS.n5356 16.0005
R7444 VSS.n5360 VSS.n5357 16.0005
R7445 VSS.n5361 VSS.n5360 16.0005
R7446 VSS.n5364 VSS.n5361 16.0005
R7447 VSS.n5366 VSS.n5364 16.0005
R7448 VSS.n5367 VSS.n5366 16.0005
R7449 VSS.n2339 VSS.n2338 16.0005
R7450 VSS.n2338 VSS.n2335 16.0005
R7451 VSS.n2335 VSS.n2334 16.0005
R7452 VSS.n2334 VSS.n2331 16.0005
R7453 VSS.n2331 VSS.n2330 16.0005
R7454 VSS.n2330 VSS.n2327 16.0005
R7455 VSS.n2327 VSS.n2326 16.0005
R7456 VSS.n2326 VSS.n2323 16.0005
R7457 VSS.n612 VSS.n611 16.0005
R7458 VSS.n611 VSS.n608 16.0005
R7459 VSS.n608 VSS.n607 16.0005
R7460 VSS.n607 VSS.n604 16.0005
R7461 VSS.n604 VSS.n603 16.0005
R7462 VSS.n603 VSS.n600 16.0005
R7463 VSS.n600 VSS.n599 16.0005
R7464 VSS.n599 VSS.n596 16.0005
R7465 VSS.n566 VSS.n564 16.0005
R7466 VSS.n564 VSS.n561 16.0005
R7467 VSS.n561 VSS.n560 16.0005
R7468 VSS.n560 VSS.n557 16.0005
R7469 VSS.n557 VSS.n556 16.0005
R7470 VSS.n556 VSS.n553 16.0005
R7471 VSS.n553 VSS.n552 16.0005
R7472 VSS.n552 VSS.n101 16.0005
R7473 VSS.n890 VSS.n888 16.0005
R7474 VSS.n888 VSS.n885 16.0005
R7475 VSS.n885 VSS.n884 16.0005
R7476 VSS.n884 VSS.n881 16.0005
R7477 VSS.n881 VSS.n880 16.0005
R7478 VSS.n880 VSS.n877 16.0005
R7479 VSS.n877 VSS.n876 16.0005
R7480 VSS.n876 VSS.n400 16.0005
R7481 VSS.n531 VSS.n530 16.0005
R7482 VSS.n530 VSS.n527 16.0005
R7483 VSS.n527 VSS.n526 16.0005
R7484 VSS.n526 VSS.n523 16.0005
R7485 VSS.n523 VSS.n522 16.0005
R7486 VSS.n522 VSS.n519 16.0005
R7487 VSS.n519 VSS.n518 16.0005
R7488 VSS.n518 VSS.n515 16.0005
R7489 VSS.n5143 VSS.n5142 16.0005
R7490 VSS.n5146 VSS.n5143 16.0005
R7491 VSS.n5147 VSS.n5146 16.0005
R7492 VSS.n5150 VSS.n5147 16.0005
R7493 VSS.n5151 VSS.n5150 16.0005
R7494 VSS.n5154 VSS.n5151 16.0005
R7495 VSS.n5156 VSS.n5154 16.0005
R7496 VSS.n5157 VSS.n5156 16.0005
R7497 VSS.n697 VSS.n696 16.0005
R7498 VSS.n696 VSS.n693 16.0005
R7499 VSS.n693 VSS.n692 16.0005
R7500 VSS.n692 VSS.n689 16.0005
R7501 VSS.n689 VSS.n688 16.0005
R7502 VSS.n688 VSS.n685 16.0005
R7503 VSS.n685 VSS.n684 16.0005
R7504 VSS.n684 VSS.n681 16.0005
R7505 VSS.n894 VSS.n893 16.0005
R7506 VSS.n897 VSS.n894 16.0005
R7507 VSS.n898 VSS.n897 16.0005
R7508 VSS.n901 VSS.n898 16.0005
R7509 VSS.n902 VSS.n901 16.0005
R7510 VSS.n905 VSS.n902 16.0005
R7511 VSS.n906 VSS.n905 16.0005
R7512 VSS.n909 VSS.n906 16.0005
R7513 VSS.n945 VSS.n942 16.0005
R7514 VSS.n946 VSS.n945 16.0005
R7515 VSS.n949 VSS.n946 16.0005
R7516 VSS.n950 VSS.n949 16.0005
R7517 VSS.n953 VSS.n950 16.0005
R7518 VSS.n954 VSS.n953 16.0005
R7519 VSS.n957 VSS.n954 16.0005
R7520 VSS.n960 VSS.n957 16.0005
R7521 VSS.n4521 VSS.n4507 16.0005
R7522 VSS.n4521 VSS.n4520 16.0005
R7523 VSS.n4520 VSS.n4519 16.0005
R7524 VSS.n4519 VSS.n4509 16.0005
R7525 VSS.n4513 VSS.n4509 16.0005
R7526 VSS.n4513 VSS.n4512 16.0005
R7527 VSS.n4512 VSS.n56 16.0005
R7528 VSS.n5480 VSS.n56 16.0005
R7529 VSS.n4314 VSS.n4313 16.0005
R7530 VSS.n4313 VSS.n4310 16.0005
R7531 VSS.n4310 VSS.n4309 16.0005
R7532 VSS.n4309 VSS.n4306 16.0005
R7533 VSS.n4306 VSS.n4305 16.0005
R7534 VSS.n4305 VSS.n4302 16.0005
R7535 VSS.n4302 VSS.n4301 16.0005
R7536 VSS.n4301 VSS.n4298 16.0005
R7537 VSS.n4394 VSS.n4393 16.0005
R7538 VSS.n4393 VSS.n4390 16.0005
R7539 VSS.n4390 VSS.n4389 16.0005
R7540 VSS.n4389 VSS.n4386 16.0005
R7541 VSS.n4386 VSS.n4385 16.0005
R7542 VSS.n4385 VSS.n4382 16.0005
R7543 VSS.n4382 VSS.n4381 16.0005
R7544 VSS.n4381 VSS.n1450 16.0005
R7545 VSS.n4582 VSS.n1409 16.0005
R7546 VSS.n1422 VSS.n1409 16.0005
R7547 VSS.n1425 VSS.n1422 16.0005
R7548 VSS.n1426 VSS.n1425 16.0005
R7549 VSS.n1429 VSS.n1426 16.0005
R7550 VSS.n1430 VSS.n1429 16.0005
R7551 VSS.n1431 VSS.n1430 16.0005
R7552 VSS.n1431 VSS.n28 16.0005
R7553 VSS.n5530 VSS.n29 16.0005
R7554 VSS.n31 VSS.n29 16.0005
R7555 VSS.n5523 VSS.n31 16.0005
R7556 VSS.n5523 VSS.n5522 16.0005
R7557 VSS.n5522 VSS.n5521 16.0005
R7558 VSS.n5521 VSS.n33 16.0005
R7559 VSS.n5516 VSS.n33 16.0005
R7560 VSS.n5516 VSS.n5515 16.0005
R7561 VSS.n3498 VSS.n1452 16.0005
R7562 VSS.n3501 VSS.n3498 16.0005
R7563 VSS.n3502 VSS.n3501 16.0005
R7564 VSS.n3505 VSS.n3502 16.0005
R7565 VSS.n3506 VSS.n3505 16.0005
R7566 VSS.n3509 VSS.n3506 16.0005
R7567 VSS.n3510 VSS.n3509 16.0005
R7568 VSS.n3511 VSS.n3510 16.0005
R7569 VSS.n3588 VSS.n3587 16.0005
R7570 VSS.n3591 VSS.n3588 16.0005
R7571 VSS.n3592 VSS.n3591 16.0005
R7572 VSS.n3595 VSS.n3592 16.0005
R7573 VSS.n3596 VSS.n3595 16.0005
R7574 VSS.n3599 VSS.n3596 16.0005
R7575 VSS.n3600 VSS.n3599 16.0005
R7576 VSS.n3603 VSS.n3600 16.0005
R7577 VSS.n3607 VSS.n3606 16.0005
R7578 VSS.n3610 VSS.n3607 16.0005
R7579 VSS.n3611 VSS.n3610 16.0005
R7580 VSS.n3614 VSS.n3611 16.0005
R7581 VSS.n3615 VSS.n3614 16.0005
R7582 VSS.n3618 VSS.n3615 16.0005
R7583 VSS.n3620 VSS.n3618 16.0005
R7584 VSS.n3621 VSS.n3620 16.0005
R7585 VSS.n3570 VSS.n1535 16.0005
R7586 VSS.n3573 VSS.n3570 16.0005
R7587 VSS.n3574 VSS.n3573 16.0005
R7588 VSS.n3577 VSS.n3574 16.0005
R7589 VSS.n3578 VSS.n3577 16.0005
R7590 VSS.n3581 VSS.n3578 16.0005
R7591 VSS.n3582 VSS.n3581 16.0005
R7592 VSS.n3585 VSS.n3582 16.0005
R7593 VSS.n1588 VSS.n1587 16.0005
R7594 VSS.n1591 VSS.n1588 16.0005
R7595 VSS.n1592 VSS.n1591 16.0005
R7596 VSS.n1595 VSS.n1592 16.0005
R7597 VSS.n1596 VSS.n1595 16.0005
R7598 VSS.n1599 VSS.n1596 16.0005
R7599 VSS.n1600 VSS.n1599 16.0005
R7600 VSS.n1603 VSS.n1600 16.0005
R7601 VSS.n1618 VSS.n1615 16.0005
R7602 VSS.n1615 VSS.n1614 16.0005
R7603 VSS.n1614 VSS.n1611 16.0005
R7604 VSS.n1611 VSS.n1610 16.0005
R7605 VSS.n1610 VSS.n1607 16.0005
R7606 VSS.n1607 VSS.n1606 16.0005
R7607 VSS.n1606 VSS.n1454 16.0005
R7608 VSS.n4500 VSS.n1454 16.0005
R7609 VSS.n3448 VSS.n3446 16.0005
R7610 VSS.n3446 VSS.n3443 16.0005
R7611 VSS.n3443 VSS.n3442 16.0005
R7612 VSS.n3442 VSS.n3439 16.0005
R7613 VSS.n3439 VSS.n3438 16.0005
R7614 VSS.n3438 VSS.n3435 16.0005
R7615 VSS.n3435 VSS.n3434 16.0005
R7616 VSS.n3434 VSS.n815 16.0005
R7617 VSS.n4810 VSS.n4809 16.0005
R7618 VSS.n4809 VSS.n4806 16.0005
R7619 VSS.n4806 VSS.n4805 16.0005
R7620 VSS.n4805 VSS.n4802 16.0005
R7621 VSS.n4802 VSS.n4801 16.0005
R7622 VSS.n4801 VSS.n4798 16.0005
R7623 VSS.n4798 VSS.n4797 16.0005
R7624 VSS.n4797 VSS.n4794 16.0005
R7625 VSS.n4890 VSS.n4889 16.0005
R7626 VSS.n4893 VSS.n4890 16.0005
R7627 VSS.n4894 VSS.n4893 16.0005
R7628 VSS.n4897 VSS.n4894 16.0005
R7629 VSS.n4898 VSS.n4897 16.0005
R7630 VSS.n4901 VSS.n4898 16.0005
R7631 VSS.n4903 VSS.n4901 16.0005
R7632 VSS.n4904 VSS.n4903 16.0005
R7633 VSS.n4828 VSS.n4827 16.0005
R7634 VSS.n4827 VSS.n4824 16.0005
R7635 VSS.n4824 VSS.n4823 16.0005
R7636 VSS.n4823 VSS.n4820 16.0005
R7637 VSS.n4820 VSS.n4819 16.0005
R7638 VSS.n4819 VSS.n4816 16.0005
R7639 VSS.n4816 VSS.n4815 16.0005
R7640 VSS.n4815 VSS.n4812 16.0005
R7641 VSS.n3753 VSS.n3752 16.0005
R7642 VSS.n3752 VSS.n3749 16.0005
R7643 VSS.n3749 VSS.n3748 16.0005
R7644 VSS.n3748 VSS.n3745 16.0005
R7645 VSS.n3745 VSS.n3744 16.0005
R7646 VSS.n3744 VSS.n3741 16.0005
R7647 VSS.n3741 VSS.n3740 16.0005
R7648 VSS.n3740 VSS.n3737 16.0005
R7649 VSS.n3704 VSS.n3701 16.0005
R7650 VSS.n3701 VSS.n3700 16.0005
R7651 VSS.n3700 VSS.n3697 16.0005
R7652 VSS.n3697 VSS.n3696 16.0005
R7653 VSS.n3696 VSS.n3693 16.0005
R7654 VSS.n3693 VSS.n3692 16.0005
R7655 VSS.n3692 VSS.n3689 16.0005
R7656 VSS.n3689 VSS.n3688 16.0005
R7657 VSS.n5303 VSS.n265 16.0005
R7658 VSS.n5303 VSS.n5302 16.0005
R7659 VSS.n5302 VSS.n5301 16.0005
R7660 VSS.n5301 VSS.n5298 16.0005
R7661 VSS.n5298 VSS.n5297 16.0005
R7662 VSS.n5297 VSS.n5294 16.0005
R7663 VSS.n5294 VSS.n5293 16.0005
R7664 VSS.n5293 VSS.n5290 16.0005
R7665 VSS.n2733 VSS.n2072 16.0005
R7666 VSS.n2733 VSS.n2732 16.0005
R7667 VSS.n2732 VSS.n2731 16.0005
R7668 VSS.n2731 VSS.n2074 16.0005
R7669 VSS.n2725 VSS.n2074 16.0005
R7670 VSS.n2725 VSS.n2724 16.0005
R7671 VSS.n2724 VSS.n2723 16.0005
R7672 VSS.n2723 VSS.n2076 16.0005
R7673 VSS.n2172 VSS.n2171 16.0005
R7674 VSS.n2173 VSS.n2172 16.0005
R7675 VSS.n2173 VSS.n2102 16.0005
R7676 VSS.n2179 VSS.n2102 16.0005
R7677 VSS.n2180 VSS.n2179 16.0005
R7678 VSS.n2181 VSS.n2180 16.0005
R7679 VSS.n2181 VSS.n2100 16.0005
R7680 VSS.n2187 VSS.n2100 16.0005
R7681 VSS.n2205 VSS.n2203 16.0005
R7682 VSS.n2203 VSS.n2200 16.0005
R7683 VSS.n2200 VSS.n2199 16.0005
R7684 VSS.n2199 VSS.n2196 16.0005
R7685 VSS.n2196 VSS.n2195 16.0005
R7686 VSS.n2195 VSS.n2192 16.0005
R7687 VSS.n2192 VSS.n2191 16.0005
R7688 VSS.n2191 VSS.n2188 16.0005
R7689 VSS.n5096 VSS.n514 16.0005
R7690 VSS.n5096 VSS.n5095 16.0005
R7691 VSS.n5095 VSS.n5094 16.0005
R7692 VSS.n5094 VSS.n5091 16.0005
R7693 VSS.n5091 VSS.n5090 16.0005
R7694 VSS.n5090 VSS.n5087 16.0005
R7695 VSS.n5087 VSS.n5086 16.0005
R7696 VSS.n5086 VSS.n5083 16.0005
R7697 VSS.n3039 VSS.n2849 16.0005
R7698 VSS.n3039 VSS.n3038 16.0005
R7699 VSS.n3038 VSS.n3037 16.0005
R7700 VSS.n3037 VSS.n2851 16.0005
R7701 VSS.n3031 VSS.n2851 16.0005
R7702 VSS.n3031 VSS.n3030 16.0005
R7703 VSS.n3030 VSS.n3029 16.0005
R7704 VSS.n3029 VSS.n2853 16.0005
R7705 VSS.n2951 VSS.n2950 16.0005
R7706 VSS.n2952 VSS.n2951 16.0005
R7707 VSS.n2952 VSS.n2881 16.0005
R7708 VSS.n2958 VSS.n2881 16.0005
R7709 VSS.n2959 VSS.n2958 16.0005
R7710 VSS.n2960 VSS.n2959 16.0005
R7711 VSS.n2960 VSS.n2879 16.0005
R7712 VSS.n2966 VSS.n2879 16.0005
R7713 VSS.n2984 VSS.n2982 16.0005
R7714 VSS.n2982 VSS.n2979 16.0005
R7715 VSS.n2979 VSS.n2978 16.0005
R7716 VSS.n2978 VSS.n2975 16.0005
R7717 VSS.n2975 VSS.n2974 16.0005
R7718 VSS.n2974 VSS.n2971 16.0005
R7719 VSS.n2971 VSS.n2970 16.0005
R7720 VSS.n2970 VSS.n2967 16.0005
R7721 VSS.n4470 VSS.n1534 16.0005
R7722 VSS.n4470 VSS.n4469 16.0005
R7723 VSS.n4469 VSS.n4468 16.0005
R7724 VSS.n4468 VSS.n4465 16.0005
R7725 VSS.n4465 VSS.n4464 16.0005
R7726 VSS.n4464 VSS.n4461 16.0005
R7727 VSS.n4461 VSS.n4460 16.0005
R7728 VSS.n4460 VSS.n4457 16.0005
R7729 VSS.n3947 VSS.n3272 16.0005
R7730 VSS.n3947 VSS.n3946 16.0005
R7731 VSS.n3946 VSS.n3945 16.0005
R7732 VSS.n3945 VSS.n3274 16.0005
R7733 VSS.n3939 VSS.n3274 16.0005
R7734 VSS.n3939 VSS.n3938 16.0005
R7735 VSS.n3938 VSS.n3937 16.0005
R7736 VSS.n3937 VSS.n3276 16.0005
R7737 VSS.n3348 VSS.n3347 16.0005
R7738 VSS.n3349 VSS.n3348 16.0005
R7739 VSS.n3349 VSS.n3304 16.0005
R7740 VSS.n3355 VSS.n3304 16.0005
R7741 VSS.n3356 VSS.n3355 16.0005
R7742 VSS.n3357 VSS.n3356 16.0005
R7743 VSS.n3357 VSS.n3302 16.0005
R7744 VSS.n3363 VSS.n3302 16.0005
R7745 VSS.n3381 VSS.n3379 16.0005
R7746 VSS.n3379 VSS.n3376 16.0005
R7747 VSS.n3376 VSS.n3375 16.0005
R7748 VSS.n3375 VSS.n3372 16.0005
R7749 VSS.n3372 VSS.n3371 16.0005
R7750 VSS.n3371 VSS.n3368 16.0005
R7751 VSS.n3368 VSS.n3367 16.0005
R7752 VSS.n3367 VSS.n3364 16.0005
R7753 VSS.n2105 VSS.n2104 16.0005
R7754 VSS.n2108 VSS.n2105 16.0005
R7755 VSS.n2109 VSS.n2108 16.0005
R7756 VSS.n2112 VSS.n2109 16.0005
R7757 VSS.n2113 VSS.n2112 16.0005
R7758 VSS.n2116 VSS.n2113 16.0005
R7759 VSS.n2117 VSS.n2116 16.0005
R7760 VSS.n2120 VSS.n2117 16.0005
R7761 VSS.n2660 VSS.n2659 16.0005
R7762 VSS.n2663 VSS.n2660 16.0005
R7763 VSS.n2664 VSS.n2663 16.0005
R7764 VSS.n2667 VSS.n2664 16.0005
R7765 VSS.n2668 VSS.n2667 16.0005
R7766 VSS.n2671 VSS.n2668 16.0005
R7767 VSS.n2673 VSS.n2671 16.0005
R7768 VSS.n2674 VSS.n2673 16.0005
R7769 VSS.n4272 VSS.n4269 16.0005
R7770 VSS.n4269 VSS.n4268 16.0005
R7771 VSS.n4268 VSS.n4265 16.0005
R7772 VSS.n4265 VSS.n4264 16.0005
R7773 VSS.n4264 VSS.n4261 16.0005
R7774 VSS.n4261 VSS.n4260 16.0005
R7775 VSS.n4260 VSS.n4257 16.0005
R7776 VSS.n4257 VSS.n1779 16.0005
R7777 VSS.n4335 VSS.n4297 16.0005
R7778 VSS.n4335 VSS.n4334 16.0005
R7779 VSS.n4334 VSS.n4333 16.0005
R7780 VSS.n4333 VSS.n4330 16.0005
R7781 VSS.n4330 VSS.n4329 16.0005
R7782 VSS.n4329 VSS.n4326 16.0005
R7783 VSS.n4326 VSS.n4325 16.0005
R7784 VSS.n4325 VSS.n4322 16.0005
R7785 VSS.n2494 VSS.n2491 16.0005
R7786 VSS.n2495 VSS.n2494 16.0005
R7787 VSS.n2498 VSS.n2495 16.0005
R7788 VSS.n2499 VSS.n2498 16.0005
R7789 VSS.n2502 VSS.n2499 16.0005
R7790 VSS.n2503 VSS.n2502 16.0005
R7791 VSS.n2506 VSS.n2503 16.0005
R7792 VSS.n2507 VSS.n2506 16.0005
R7793 VSS.n2408 VSS.n2405 16.0005
R7794 VSS.n2405 VSS.n2404 16.0005
R7795 VSS.n2404 VSS.n2401 16.0005
R7796 VSS.n2401 VSS.n2400 16.0005
R7797 VSS.n2400 VSS.n2397 16.0005
R7798 VSS.n2397 VSS.n2396 16.0005
R7799 VSS.n2396 VSS.n2393 16.0005
R7800 VSS.n2393 VSS.n1408 16.0005
R7801 VSS.n1873 VSS.n1872 13.7392
R7802 VSS.n5352 VSS.n168 13.6894
R7803 VSS.n680 VSS.n531 13.6894
R7804 VSS.n5142 VSS.n422 13.6894
R7805 VSS.n4507 VSS.n4506 13.6894
R7806 VSS.n4394 VSS.n1689 13.6894
R7807 VSS.n3587 VSS.n3586 13.6894
R7808 VSS.n3606 VSS.n3604 13.6894
R7809 VSS.n4811 VSS.n4810 13.6894
R7810 VSS.n4889 VSS.n837 13.6894
R7811 VSS.n4094 VSS.n4081 13.5116
R7812 VSS.n3251 VSS.n1953 13.5116
R7813 VSS.n3111 VSS.n3109 13.5116
R7814 VSS.n2828 VSS.n2029 13.5116
R7815 VSS.n2659 VSS.n2584 13.5116
R7816 VSS.n4793 VSS.n4792 13.3338
R7817 VSS.n4768 VSS.n1128 13.3338
R7818 VSS.n5289 VSS.n266 13.3338
R7819 VSS.n5082 VSS.n697 13.3338
R7820 VSS.n4321 VSS.n4314 13.3338
R7821 VSS.n4456 VSS.n1535 13.3338
R7822 VSS.n4829 VSS.n4828 13.3338
R7823 VSS.n2711 VSS.n265 13.3338
R7824 VSS.n2675 VSS.n2072 13.3338
R7825 VSS.n3017 VSS.n514 13.3338
R7826 VSS.n2849 VSS.n2848 13.3338
R7827 VSS.n3925 VSS.n1534 13.3338
R7828 VSS.n3272 VSS.n3271 13.3338
R7829 VSS.n4273 VSS.n4272 13.3338
R7830 VSS.n4297 VSS.n4296 13.3338
R7831 VSS.n4632 VSS.n4631 12.1065
R7832 VSS.n4673 VSS.n4672 11.6369
R7833 VSS.n4672 VSS.n4671 11.6369
R7834 VSS.n4671 VSS.n1365 11.6369
R7835 VSS.n1367 VSS.n1365 11.6369
R7836 VSS.n2522 VSS.n1367 11.6369
R7837 VSS.n2523 VSS.n2522 11.6369
R7838 VSS.n2523 VSS.n2518 11.6369
R7839 VSS.n2530 VSS.n2518 11.6369
R7840 VSS.n2259 VSS.n2256 11.6369
R7841 VSS.n2380 VSS.n2259 11.6369
R7842 VSS.n2380 VSS.n2379 11.6369
R7843 VSS.n2379 VSS.n2378 11.6369
R7844 VSS.n2378 VSS.n2260 11.6369
R7845 VSS.n2372 VSS.n2260 11.6369
R7846 VSS.n2372 VSS.n2371 11.6369
R7847 VSS.n2371 VSS.n2370 11.6369
R7848 VSS.n2291 VSS.n2289 11.6369
R7849 VSS.n2291 VSS.n2290 11.6369
R7850 VSS.n2290 VSS.n162 11.6369
R7851 VSS.n5383 VSS.n162 11.6369
R7852 VSS.n5383 VSS.n5382 11.6369
R7853 VSS.n5382 VSS.n5381 11.6369
R7854 VSS.n5381 VSS.n163 11.6369
R7855 VSS.n5375 VSS.n163 11.6369
R7856 VSS.n2322 VSS.n2266 11.6369
R7857 VSS.n2316 VSS.n2266 11.6369
R7858 VSS.n2316 VSS.n2315 11.6369
R7859 VSS.n2315 VSS.n2314 11.6369
R7860 VSS.n2314 VSS.n2273 11.6369
R7861 VSS.n2308 VSS.n2273 11.6369
R7862 VSS.n2308 VSS.n2307 11.6369
R7863 VSS.n2307 VSS.n2306 11.6369
R7864 VSS.n2685 VSS.n2577 11.6369
R7865 VSS.n2691 VSS.n2577 11.6369
R7866 VSS.n2692 VSS.n2691 11.6369
R7867 VSS.n2693 VSS.n2692 11.6369
R7868 VSS.n2693 VSS.n2575 11.6369
R7869 VSS.n2699 VSS.n2575 11.6369
R7870 VSS.n2700 VSS.n2699 11.6369
R7871 VSS.n2702 VSS.n2700 11.6369
R7872 VSS.n2565 VSS.n2564 11.6369
R7873 VSS.n2564 VSS.n2563 11.6369
R7874 VSS.n2563 VSS.n2245 11.6369
R7875 VSS.n2247 VSS.n2245 11.6369
R7876 VSS.n2250 VSS.n2247 11.6369
R7877 VSS.n2553 VSS.n2250 11.6369
R7878 VSS.n2553 VSS.n2552 11.6369
R7879 VSS.n2552 VSS.n2551 11.6369
R7880 VSS.n2615 VSS.n2591 11.6369
R7881 VSS.n2615 VSS.n2614 11.6369
R7882 VSS.n2614 VSS.n2613 11.6369
R7883 VSS.n2613 VSS.n2595 11.6369
R7884 VSS.n2603 VSS.n2595 11.6369
R7885 VSS.n2605 VSS.n2603 11.6369
R7886 VSS.n2605 VSS.n2604 11.6369
R7887 VSS.n2604 VSS.n2581 11.6369
R7888 VSS.n4161 VSS.n4160 11.6369
R7889 VSS.n4161 VSS.n1864 11.6369
R7890 VSS.n4167 VSS.n1864 11.6369
R7891 VSS.n4168 VSS.n4167 11.6369
R7892 VSS.n4170 VSS.n4168 11.6369
R7893 VSS.n4170 VSS.n4169 11.6369
R7894 VSS.n4169 VSS.n1861 11.6369
R7895 VSS.n1861 VSS.n1853 11.6369
R7896 VSS.n4210 VSS.n1854 11.6369
R7897 VSS.n4204 VSS.n1854 11.6369
R7898 VSS.n4204 VSS.n4203 11.6369
R7899 VSS.n4203 VSS.n4202 11.6369
R7900 VSS.n4202 VSS.n4185 11.6369
R7901 VSS.n4189 VSS.n4185 11.6369
R7902 VSS.n4195 VSS.n4189 11.6369
R7903 VSS.n4195 VSS.n4194 11.6369
R7904 VSS.n2534 VSS.n2532 11.6369
R7905 VSS.n2535 VSS.n2534 11.6369
R7906 VSS.n2535 VSS.n1382 11.6369
R7907 VSS.n4654 VSS.n1382 11.6369
R7908 VSS.n4654 VSS.n4653 11.6369
R7909 VSS.n4653 VSS.n4652 11.6369
R7910 VSS.n4652 VSS.n1383 11.6369
R7911 VSS.n4646 VSS.n1383 11.6369
R7912 VSS.n4589 VSS.n4588 11.6369
R7913 VSS.n4614 VSS.n4589 11.6369
R7914 VSS.n4614 VSS.n4613 11.6369
R7915 VSS.n4613 VSS.n4612 11.6369
R7916 VSS.n4612 VSS.n4590 11.6369
R7917 VSS.n4594 VSS.n4590 11.6369
R7918 VSS.n4604 VSS.n4594 11.6369
R7919 VSS.n4604 VSS.n4603 11.6369
R7920 VSS.n4603 VSS.n4602 11.6369
R7921 VSS.n5544 VSS.n5543 11.6369
R7922 VSS.n5545 VSS.n5544 11.6369
R7923 VSS.n5545 VSS.n11 11.6369
R7924 VSS.n5551 VSS.n11 11.6369
R7925 VSS.n5552 VSS.n5551 11.6369
R7926 VSS.n5554 VSS.n5552 11.6369
R7927 VSS.n5554 VSS.n5553 11.6369
R7928 VSS.n5553 VSS.n8 11.6369
R7929 VSS.n4986 VSS.n765 11.5043
R7930 VSS.n1684 VSS.n1654 11.5043
R7931 VSS.n675 VSS.n645 11.5043
R7932 VSS.n5543 VSS.n18 11.0106
R7933 VSS.n4673 VSS.n1361 10.9261
R7934 VSS.n4602 VSS.n4596 10.9063
R7935 VSS.n2565 VSS.n2244 10.8998
R7936 VSS.t14 VSS.t81 10.8468
R7937 VSS.t16 VSS.t3 10.8468
R7938 VSS.n638 VSS.n612 10.3116
R7939 VSS.n595 VSS.n566 10.3116
R7940 VSS.n961 VSS.n890 10.3116
R7941 VSS.n942 VSS.n941 10.3116
R7942 VSS.n4583 VSS.n4582 10.3116
R7943 VSS.n5531 VSS.n5530 10.3116
R7944 VSS.n4501 VSS.n1452 10.3116
R7945 VSS.n1650 VSS.n1618 10.3116
R7946 VSS.n3449 VSS.n3448 10.3116
R7947 VSS.n3736 VSS.n3704 10.3116
R7948 VSS.n4148 VSS.n4147 10.1338
R7949 VSS.n3221 VSS.n3219 10.1338
R7950 VSS.n1979 VSS.n1978 10.1338
R7951 VSS.n2883 VSS.n1995 10.1338
R7952 VSS.n2104 VSS.n2038 10.1338
R7953 VSS.n2289 VSS.n2277 10.0853
R7954 VSS.n2622 VSS.n2591 10.0103
R7955 VSS.n4160 VSS.n4159 10.0103
R7956 VSS.n2436 VSS.n1849 9.95606
R7957 VSS.n3416 VSS.n1153 9.95606
R7958 VSS.n3866 VSS.n3829 9.95606
R7959 VSS.n534 VSS.n291 9.95606
R7960 VSS.n893 VSS.n719 9.95606
R7961 VSS.n1587 VSS.n1556 9.95606
R7962 VSS.n3811 VSS.n3753 9.95606
R7963 VSS.n2171 VSS.n2121 9.95606
R7964 VSS.n2206 VSS.n2205 9.95606
R7965 VSS.n2950 VSS.n2900 9.95606
R7966 VSS.n2985 VSS.n2984 9.95606
R7967 VSS.n3347 VSS.n1922 9.95606
R7968 VSS.n3382 VSS.n3381 9.95606
R7969 VSS.n2491 VSS.n2490 9.95606
R7970 VSS.n2409 VSS.n2408 9.95606
R7971 VSS.n2256 VSS.n2251 9.82676
R7972 VSS.n2685 VSS.n2684 9.82676
R7973 VSS.n4211 VSS.n4210 9.82676
R7974 VSS.n2532 VSS.n2531 9.82676
R7975 VSS.n4588 VSS.n4586 9.7416
R7976 VSS.n4622 VSS.n1398 9.32831
R7977 VSS.n1885 VSS.t23 8.7005
R7978 VSS.n1885 VSS.t77 8.7005
R7979 VSS.n1884 VSS.t25 8.7005
R7980 VSS.n1884 VSS.t21 8.7005
R7981 VSS.n4194 VSS.n4193 8.13406
R7982 VSS.n2702 VSS.n2701 8.00427
R7983 VSS.n4646 VSS.n4645 7.95163
R7984 VSS.n2490 VSS.n2452 7.11161
R7985 VSS.n3866 VSS.n3432 7.11161
R7986 VSS.n638 VSS.n550 7.11161
R7987 VSS.n596 VSS.n595 7.11161
R7988 VSS.n5419 VSS.n101 7.11161
R7989 VSS.n5206 VSS.n400 7.11161
R7990 VSS.n941 VSS.n909 7.11161
R7991 VSS.n961 VSS.n960 7.11161
R7992 VSS.n5531 VSS.n28 7.11161
R7993 VSS.n5515 VSS.n5514 7.11161
R7994 VSS.n3511 VSS.n62 7.11161
R7995 VSS.n1650 VSS.n1603 7.11161
R7996 VSS.n4501 VSS.n4500 7.11161
R7997 VSS.n4953 VSS.n815 7.11161
R7998 VSS.n3737 VSS.n3736 7.11161
R7999 VSS.n3688 VSS.n3449 7.11161
R8000 VSS.n2206 VSS.n2187 7.11161
R8001 VSS.n2985 VSS.n2966 7.11161
R8002 VSS.n3382 VSS.n3363 7.11161
R8003 VSS.n4583 VSS.n1408 7.11161
R8004 VSS.n4193 VSS.n4190 7.06798
R8005 VSS.n4679 VSS.n1361 7.06798
R8006 VSS.n1897 VSS.n1871 7.02795
R8007 VSS.n4596 VSS.n4595 6.94026
R8008 VSS.n5537 VSS.n18 6.94026
R8009 VSS.n4130 VSS.n1849 6.93383
R8010 VSS.n3203 VSS.n1922 6.93383
R8011 VSS.n1961 VSS.n1153 6.93383
R8012 VSS.n2900 VSS.n2899 6.93383
R8013 VSS.n3812 VSS.n3811 6.93383
R8014 VSS.n2188 VSS.n291 6.93383
R8015 VSS.n2967 VSS.n719 6.93383
R8016 VSS.n3364 VSS.n1556 6.93383
R8017 VSS.n2121 VSS.n2120 6.93383
R8018 VSS.n2507 VSS.n2409 6.93383
R8019 VSS.n2701 VSS.n2572 6.8987
R8020 VSS.n2244 VSS.n2240 6.8987
R8021 VSS.n4645 VSS.n4644 6.8987
R8022 VSS.n4680 VSS.n4679 6.59682
R8023 VSS.n5537 VSS.n5536 6.47761
R8024 VSS.n2709 VSS.n2240 6.43882
R8025 VSS.n4586 VSS.n4585 6.43882
R8026 VSS.n4585 VSS.n4584 6.28553
R8027 VSS.n24 VSS.n22 6.16917
R8028 VSS VSS.n4630 6.09612
R8029 VSS.n4068 VSS.n4067 5.81868
R8030 VSS.n4067 VSS.n4066 5.81868
R8031 VSS.n4066 VSS.n4003 5.81868
R8032 VSS.n4061 VSS.n4003 5.81868
R8033 VSS.n4061 VSS.n4060 5.81868
R8034 VSS.n4060 VSS.n4059 5.81868
R8035 VSS.n4059 VSS.n4005 5.81868
R8036 VSS.n4053 VSS.n4005 5.81868
R8037 VSS.n5248 VSS.n5247 5.81868
R8038 VSS.n5247 VSS.n5245 5.81868
R8039 VSS.n5245 VSS.n309 5.81868
R8040 VSS.n313 VSS.n309 5.81868
R8041 VSS.n315 VSS.n313 5.81868
R8042 VSS.n317 VSS.n315 5.81868
R8043 VSS.n319 VSS.n317 5.81868
R8044 VSS.n5238 VSS.n319 5.81868
R8045 VSS.n4415 VSS.n4414 5.81868
R8046 VSS.n4414 VSS.n4412 5.81868
R8047 VSS.n4412 VSS.n1573 5.81868
R8048 VSS.n1577 VSS.n1573 5.81868
R8049 VSS.n1579 VSS.n1577 5.81868
R8050 VSS.n1581 VSS.n1579 5.81868
R8051 VSS.n1583 VSS.n1581 5.81868
R8052 VSS.n4405 VSS.n1583 5.81868
R8053 VSS.n1681 VSS.n1652 5.81868
R8054 VSS.n1681 VSS.n1680 5.81868
R8055 VSS.n1680 VSS.n1679 5.81868
R8056 VSS.n1679 VSS.n1657 5.81868
R8057 VSS.n1659 VSS.n1657 5.81868
R8058 VSS.n1662 VSS.n1659 5.81868
R8059 VSS.n1669 VSS.n1662 5.81868
R8060 VSS.n1669 VSS.n1668 5.81868
R8061 VSS.n1668 VSS.n1667 5.81868
R8062 VSS.n5446 VSS.n5445 5.81868
R8063 VSS.n5450 VSS.n5446 5.81868
R8064 VSS.n5451 VSS.n5450 5.81868
R8065 VSS.n5455 VSS.n5451 5.81868
R8066 VSS.n5457 VSS.n5455 5.81868
R8067 VSS.n5458 VSS.n5457 5.81868
R8068 VSS.n5458 VSS.n63 5.81868
R8069 VSS.n5466 VSS.n63 5.81868
R8070 VSS.n5004 VSS.n5003 5.81868
R8071 VSS.n5003 VSS.n5001 5.81868
R8072 VSS.n5001 VSS.n749 5.81868
R8073 VSS.n753 VSS.n749 5.81868
R8074 VSS.n755 VSS.n753 5.81868
R8075 VSS.n757 VSS.n755 5.81868
R8076 VSS.n759 VSS.n757 5.81868
R8077 VSS.n4994 VSS.n759 5.81868
R8078 VSS.n4983 VSS.n763 5.81868
R8079 VSS.n4983 VSS.n4982 5.81868
R8080 VSS.n4982 VSS.n4981 5.81868
R8081 VSS.n4981 VSS.n768 5.81868
R8082 VSS.n770 VSS.n768 5.81868
R8083 VSS.n773 VSS.n770 5.81868
R8084 VSS.n4971 VSS.n773 5.81868
R8085 VSS.n4971 VSS.n4970 5.81868
R8086 VSS.n4970 VSS.n4969 5.81868
R8087 VSS.n5041 VSS.n5040 5.81868
R8088 VSS.n5040 VSS.n5038 5.81868
R8089 VSS.n5038 VSS.n5020 5.81868
R8090 VSS.n5024 VSS.n5020 5.81868
R8091 VSS.n5026 VSS.n5024 5.81868
R8092 VSS.n5028 VSS.n5026 5.81868
R8093 VSS.n5030 VSS.n5028 5.81868
R8094 VSS.n5031 VSS.n5030 5.81868
R8095 VSS.n5227 VSS.n335 5.81868
R8096 VSS.n348 VSS.n335 5.81868
R8097 VSS.n350 VSS.n348 5.81868
R8098 VSS.n352 VSS.n350 5.81868
R8099 VSS.n353 VSS.n352 5.81868
R8100 VSS.n355 VSS.n353 5.81868
R8101 VSS.n355 VSS.n354 5.81868
R8102 VSS.n354 VSS.n343 5.81868
R8103 VSS.n5220 VSS.n343 5.81868
R8104 VSS.n379 VSS.n377 5.81868
R8105 VSS.n381 VSS.n379 5.81868
R8106 VSS.n383 VSS.n381 5.81868
R8107 VSS.n384 VSS.n383 5.81868
R8108 VSS.n385 VSS.n384 5.81868
R8109 VSS.n385 VSS.n369 5.81868
R8110 VSS.n391 VSS.n369 5.81868
R8111 VSS.n393 VSS.n391 5.81868
R8112 VSS.n794 VSS.n792 5.81868
R8113 VSS.n796 VSS.n794 5.81868
R8114 VSS.n798 VSS.n796 5.81868
R8115 VSS.n799 VSS.n798 5.81868
R8116 VSS.n800 VSS.n799 5.81868
R8117 VSS.n800 VSS.n784 5.81868
R8118 VSS.n806 VSS.n784 5.81868
R8119 VSS.n808 VSS.n806 5.81868
R8120 VSS.n142 VSS.n140 5.81868
R8121 VSS.n144 VSS.n142 5.81868
R8122 VSS.n146 VSS.n144 5.81868
R8123 VSS.n148 VSS.n146 5.81868
R8124 VSS.n150 VSS.n148 5.81868
R8125 VSS.n151 VSS.n150 5.81868
R8126 VSS.n154 VSS.n151 5.81868
R8127 VSS.n154 VSS.n153 5.81868
R8128 VSS.n672 VSS.n644 5.81868
R8129 VSS.n672 VSS.n671 5.81868
R8130 VSS.n671 VSS.n670 5.81868
R8131 VSS.n670 VSS.n648 5.81868
R8132 VSS.n650 VSS.n648 5.81868
R8133 VSS.n653 VSS.n650 5.81868
R8134 VSS.n660 VSS.n653 5.81868
R8135 VSS.n660 VSS.n659 5.81868
R8136 VSS.n659 VSS.n658 5.81868
R8137 VSS.n4703 VSS.n1206 5.81868
R8138 VSS.n4703 VSS.n4702 5.81868
R8139 VSS.n4702 VSS.n4701 5.81868
R8140 VSS.n4701 VSS.n1213 5.81868
R8141 VSS.n1215 VSS.n1213 5.81868
R8142 VSS.n1218 VSS.n1215 5.81868
R8143 VSS.n4693 VSS.n1218 5.81868
R8144 VSS.n4693 VSS.n4692 5.81868
R8145 VSS.n1229 VSS.n1225 5.81868
R8146 VSS.n1249 VSS.n1229 5.81868
R8147 VSS.n1249 VSS.n1248 5.81868
R8148 VSS.n1248 VSS.n1231 5.81868
R8149 VSS.n1232 VSS.n1231 5.81868
R8150 VSS.n1240 VSS.n1232 5.81868
R8151 VSS.n1240 VSS.n1239 5.81868
R8152 VSS.n1239 VSS.n1234 5.81868
R8153 VSS.n1283 VSS.n1279 5.81868
R8154 VSS.n1284 VSS.n1283 5.81868
R8155 VSS.n1288 VSS.n1284 5.81868
R8156 VSS.n1289 VSS.n1288 5.81868
R8157 VSS.n1293 VSS.n1289 5.81868
R8158 VSS.n1294 VSS.n1293 5.81868
R8159 VSS.n1298 VSS.n1294 5.81868
R8160 VSS.n1301 VSS.n1298 5.81868
R8161 VSS.n1331 VSS.n1308 5.81868
R8162 VSS.n1331 VSS.n1330 5.81868
R8163 VSS.n1330 VSS.n1310 5.81868
R8164 VSS.n1311 VSS.n1310 5.81868
R8165 VSS.n1322 VSS.n1311 5.81868
R8166 VSS.n1322 VSS.n1321 5.81868
R8167 VSS.n1321 VSS.n1313 5.81868
R8168 VSS.n1314 VSS.n1313 5.81868
R8169 VSS.n4036 VSS.n4029 5.81868
R8170 VSS.n4036 VSS.n4035 5.81868
R8171 VSS.n4035 VSS.n4033 5.81868
R8172 VSS.n4033 VSS.n4031 5.81868
R8173 VSS.n4031 VSS.n4022 5.81868
R8174 VSS.n4042 VSS.n4022 5.81868
R8175 VSS.n4043 VSS.n4042 5.81868
R8176 VSS.n4044 VSS.n4043 5.81868
R8177 VSS.n4724 VSS.n1161 5.81868
R8178 VSS.n4724 VSS.n4723 5.81868
R8179 VSS.n4723 VSS.n4722 5.81868
R8180 VSS.n4722 VSS.n1169 5.81868
R8181 VSS.n3909 VSS.n1169 5.81868
R8182 VSS.n3911 VSS.n3909 5.81868
R8183 VSS.n3911 VSS.n3910 5.81868
R8184 VSS.n3910 VSS.n3905 5.81868
R8185 VSS.n3899 VSS.n3873 5.81868
R8186 VSS.n3874 VSS.n3873 5.81868
R8187 VSS.n3891 VSS.n3874 5.81868
R8188 VSS.n3891 VSS.n3890 5.81868
R8189 VSS.n3890 VSS.n3876 5.81868
R8190 VSS.n3877 VSS.n3876 5.81868
R8191 VSS.n3882 VSS.n3877 5.81868
R8192 VSS.n3882 VSS.n3881 5.81868
R8193 VSS.n3983 VSS.n3981 5.81868
R8194 VSS.n3985 VSS.n3983 5.81868
R8195 VSS.n3987 VSS.n3985 5.81868
R8196 VSS.n3988 VSS.n3987 5.81868
R8197 VSS.n3989 VSS.n3988 5.81868
R8198 VSS.n3989 VSS.n3974 5.81868
R8199 VSS.n3995 VSS.n3974 5.81868
R8200 VSS.n3997 VSS.n3995 5.81868
R8201 VSS.n3079 VSS.n3077 5.81868
R8202 VSS.n3081 VSS.n3079 5.81868
R8203 VSS.n3083 VSS.n3081 5.81868
R8204 VSS.n3084 VSS.n3083 5.81868
R8205 VSS.n3084 VSS.n3073 5.81868
R8206 VSS.n3091 VSS.n3073 5.81868
R8207 VSS.n3092 VSS.n3091 5.81868
R8208 VSS.n3093 VSS.n3092 5.81868
R8209 VSS.n3164 VSS.n3162 5.81868
R8210 VSS.n3166 VSS.n3164 5.81868
R8211 VSS.n3168 VSS.n3166 5.81868
R8212 VSS.n3170 VSS.n3168 5.81868
R8213 VSS.n3172 VSS.n3170 5.81868
R8214 VSS.n3174 VSS.n3172 5.81868
R8215 VSS.n3174 VSS.n3173 5.81868
R8216 VSS.n3173 VSS.n1162 5.81868
R8217 VSS.n2785 VSS.n2784 5.81868
R8218 VSS.n2784 VSS.n2783 5.81868
R8219 VSS.n2783 VSS.n2763 5.81868
R8220 VSS.n2765 VSS.n2763 5.81868
R8221 VSS.n2771 VSS.n2765 5.81868
R8222 VSS.n2773 VSS.n2771 5.81868
R8223 VSS.n2773 VSS.n2772 5.81868
R8224 VSS.n2772 VSS.n1207 5.81868
R8225 VSS.n5445 VSS.n5441 5.51409
R8226 VSS.n377 VSS.n375 5.51409
R8227 VSS.n792 VSS.n790 5.51409
R8228 VSS.n140 VSS.n85 5.51409
R8229 VSS.n5421 VSS.n5420 5.50178
R8230 VSS.n5208 VSS.n5207 5.50178
R8231 VSS.n4955 VSS.n4954 5.50178
R8232 VSS.n5469 VSS.n5468 5.50178
R8233 VSS.n5513 VSS.n6 5.50178
R8234 VSS.n2759 VSS.n2758 5.47847
R8235 VSS.n3065 VSS.n3064 5.47847
R8236 VSS.n3151 VSS.n3150 5.47847
R8237 VSS.n3220 VSS.n1913 5.47847
R8238 VSS.n4159 VSS.n1868 5.47847
R8239 VSS.n1667 VSS.n1663 5.46332
R8240 VSS.n4969 VSS.n774 5.46332
R8241 VSS.n5220 VSS.n5219 5.46332
R8242 VSS.n658 VSS.n82 5.46332
R8243 VSS.n1257 VSS.n1225 5.46332
R8244 VSS.n1308 VSS.n1278 5.46332
R8245 VSS.n4029 VSS.n4028 5.46332
R8246 VSS.n3900 VSS.n3899 5.46332
R8247 VSS.n5374 VSS.n5373 5.22944
R8248 VSS.n5426 VSS.n96 5.22944
R8249 VSS.n5213 VSS.n395 5.22944
R8250 VSS.n4960 VSS.n810 5.22944
R8251 VSS.n5477 VSS.n57 5.22944
R8252 VSS.n2623 VSS.n2622 5.20728
R8253 VSS.n2792 VSS.n2791 5.20728
R8254 VSS.n3112 VSS.n3098 5.20728
R8255 VSS.n3184 VSS.n3183 5.20728
R8256 VSS.n4080 VSS.n1911 5.20728
R8257 VSS.n3981 VSS.n3979 4.97828
R8258 VSS.n3077 VSS.n1993 4.97828
R8259 VSS.n3162 VSS.n1959 4.97828
R8260 VSS.n2785 VSS.n2036 4.97828
R8261 VSS.n4068 VSS.n3998 4.91363
R8262 VSS.n5248 VSS.n299 4.91363
R8263 VSS.n4415 VSS.n1563 4.91363
R8264 VSS.n5004 VSS.n740 4.91363
R8265 VSS.n5041 VSS.n727 4.91363
R8266 VSS.n4710 VSS.n1206 4.91363
R8267 VSS.n1279 VSS.n1196 4.91363
R8268 VSS.n4731 VSS.n1161 4.91363
R8269 VSS.n1686 VSS.n1652 4.90491
R8270 VSS.n4988 VSS.n763 4.90491
R8271 VSS.n5228 VSS.n5227 4.90491
R8272 VSS.n677 VSS.n644 4.90491
R8273 VSS.n1360 VSS.n1357 4.24099
R8274 VSS.n2710 VSS.n2239 4.13942
R8275 VSS.n4053 VSS.n4052 4.06728
R8276 VSS.n4692 VSS.n4691 4.06728
R8277 VSS.n1302 VSS.n1301 4.06728
R8278 VSS.n3918 VSS.n3905 4.06728
R8279 VSS.n5238 VSS.n5237 4.0419
R8280 VSS.n4405 VSS.n4404 4.0419
R8281 VSS.n4994 VSS.n4993 4.0419
R8282 VSS.n5031 VSS.n331 4.0419
R8283 VSS.n5412 VSS.n123 4.03114
R8284 VSS.n5411 VSS.n124 4.03114
R8285 VSS.n132 VSS.n130 4.03114
R8286 VSS.n5405 VSS.n5404 4.03114
R8287 VSS.n5401 VSS.n133 4.03114
R8288 VSS.n5392 VSS.n5388 4.03114
R8289 VSS.n5394 VSS.n5393 4.03114
R8290 VSS.n5417 VSS.n102 4.03114
R8291 VSS.n5199 VSS.n5159 4.03114
R8292 VSS.n5198 VSS.n5160 4.03114
R8293 VSS.n5170 VSS.n5168 4.03114
R8294 VSS.n5192 VSS.n5191 4.03114
R8295 VSS.n5188 VSS.n5171 4.03114
R8296 VSS.n5179 VSS.n5175 4.03114
R8297 VSS.n5181 VSS.n5180 4.03114
R8298 VSS.n5204 VSS.n401 4.03114
R8299 VSS.n4946 VSS.n4906 4.03114
R8300 VSS.n4945 VSS.n4907 4.03114
R8301 VSS.n4917 VSS.n4915 4.03114
R8302 VSS.n4939 VSS.n4938 4.03114
R8303 VSS.n4935 VSS.n4918 4.03114
R8304 VSS.n4926 VSS.n4922 4.03114
R8305 VSS.n4928 VSS.n4927 4.03114
R8306 VSS.n4951 VSS.n816 4.03114
R8307 VSS.n3668 VSS.n3623 4.03114
R8308 VSS.n3667 VSS.n3624 4.03114
R8309 VSS.n3634 VSS.n3632 4.03114
R8310 VSS.n3661 VSS.n3660 4.03114
R8311 VSS.n3657 VSS.n3635 4.03114
R8312 VSS.n3643 VSS.n3639 4.03114
R8313 VSS.n3650 VSS.n3649 4.03114
R8314 VSS.n3646 VSS.n3644 4.03114
R8315 VSS.n5478 VSS.n53 4.03114
R8316 VSS.n5489 VSS.n5488 4.03114
R8317 VSS.n5485 VSS.n54 4.03114
R8318 VSS.n50 VSS.n49 4.03114
R8319 VSS.n5498 VSS.n47 4.03114
R8320 VSS.n44 VSS.n40 4.03114
R8321 VSS.n5506 VSS.n5505 4.03114
R8322 VSS.n41 VSS.n36 4.03114
R8323 VSS.n5389 VSS 3.97667
R8324 VSS.n5176 VSS 3.97667
R8325 VSS.n4923 VSS 3.97667
R8326 VSS.n3640 VSS 3.97667
R8327 VSS VSS.n45 3.97667
R8328 VSS.n4792 VSS.n1055 3.73383
R8329 VSS.n2356 VSS.n2355 3.73383
R8330 VSS.n5368 VSS.n5367 3.73383
R8331 VSS.n2323 VSS.n168 3.73383
R8332 VSS.n515 VSS.n422 3.73383
R8333 VSS.n5158 VSS.n5157 3.73383
R8334 VSS.n681 VSS.n680 3.73383
R8335 VSS.n5480 VSS.n5479 3.73383
R8336 VSS.n4298 VSS.n1689 3.73383
R8337 VSS.n4506 VSS.n1450 3.73383
R8338 VSS.n3604 VSS.n3603 3.73383
R8339 VSS.n3622 VSS.n3621 3.73383
R8340 VSS.n3586 VSS.n3585 3.73383
R8341 VSS.n4794 VSS.n837 3.73383
R8342 VSS.n4905 VSS.n4904 3.73383
R8343 VSS.n4812 VSS.n4811 3.73383
R8344 VSS.n2711 VSS.n2076 3.73383
R8345 VSS.n3017 VSS.n2853 3.73383
R8346 VSS.n3925 VSS.n3276 3.73383
R8347 VSS.n4296 VSS.n1779 3.73383
R8348 VSS VSS.n5566 3.70844
R8349 VSS.n4680 VSS.n1360 3.6913
R8350 VSS VSS.n2 3.67867
R8351 VSS.n2710 VSS.n2709 3.6029
R8352 VSS.n4274 VSS.n4273 3.55606
R8353 VSS.n3271 VSS.n3266 3.55606
R8354 VSS.n4770 VSS.n4768 3.55606
R8355 VSS.n2848 VSS.n2843 3.55606
R8356 VSS.n4830 VSS.n4829 3.55606
R8357 VSS.n5290 VSS.n5289 3.55606
R8358 VSS.n5083 VSS.n5082 3.55606
R8359 VSS.n4457 VSS.n4456 3.55606
R8360 VSS.n2675 VSS.n2674 3.55606
R8361 VSS.n4322 VSS.n4321 3.55606
R8362 VSS.n4404 VSS.n4403 3.53424
R8363 VSS.n1663 VSS.n74 3.53424
R8364 VSS.n5441 VSS.n5440 3.53424
R8365 VSS.n4993 VSS.n4992 3.53424
R8366 VSS.n5232 VSS.n331 3.53424
R8367 VSS.n5219 VSS.n359 3.53424
R8368 VSS.n375 VSS.n361 3.53424
R8369 VSS.n3476 VSS.n774 3.53424
R8370 VSS.n790 VSS.n776 3.53424
R8371 VSS.n5434 VSS.n82 3.53424
R8372 VSS.n5430 VSS.n85 3.53424
R8373 VSS.n5237 VSS.n5236 3.53424
R8374 VSS.n4691 VSS.n1219 3.53424
R8375 VSS.n1258 VSS.n1257 3.53424
R8376 VSS.n1303 VSS.n1302 3.53424
R8377 VSS.n1339 VSS.n1278 3.53424
R8378 VSS.n4052 VSS.n4051 3.53424
R8379 VSS.n4028 VSS.n4015 3.53424
R8380 VSS.n3920 VSS.n3918 3.53424
R8381 VSS.n3900 VSS.n3869 3.53424
R8382 VSS.n1687 VSS.n1686 3.29866
R8383 VSS.n5440 VSS.n70 3.29866
R8384 VSS.n4989 VSS.n4988 3.29866
R8385 VSS.n5229 VSS.n5228 3.29866
R8386 VSS.n966 VSS.n361 3.29866
R8387 VSS.n3680 VSS.n776 3.29866
R8388 VSS.n5431 VSS.n5430 3.29866
R8389 VSS.n678 VSS.n677 3.29866
R8390 VSS.n4686 VSS.n1258 3.29866
R8391 VSS.n1340 VSS.n1339 3.29866
R8392 VSS.n4015 VSS.n4014 3.29866
R8393 VSS.n3923 VSS.n3869 3.29866
R8394 VSS.n2546 VSS.n1 3.22364
R8395 VSS.n1687 VSS.n1651 3.22013
R8396 VSS.n4989 VSS.n761 3.22013
R8397 VSS.n5229 VSS.n332 3.22013
R8398 VSS.n679 VSS.n678 3.22013
R8399 VSS.n4623 VSS.n4622 3.15497
R8400 VSS.n4502 VSS.n1451 3.1416
R8401 VSS.n847 VSS.n846 3.1416
R8402 VSS.n3478 VSS.n3477 3.1416
R8403 VSS.n5433 VSS.n83 3.1416
R8404 VSS.n4630 VSS.n4629 3.1005
R8405 VSS.n5373 VSS.n5368 2.83284
R8406 VSS.n5158 VSS.n96 2.83284
R8407 VSS.n4905 VSS.n395 2.83284
R8408 VSS.n3622 VSS.n810 2.83284
R8409 VSS.n5479 VSS.n5477 2.83284
R8410 VSS.n2623 VSS.n2584 2.82084
R8411 VSS.n2792 VSS.n2029 2.82084
R8412 VSS.n3112 VSS.n3111 2.82084
R8413 VSS.n3184 VSS.n1953 2.82084
R8414 VSS.n4081 VSS.n4080 2.82084
R8415 VSS.n5426 VSS.n95 2.77837
R8416 VSS.n5213 VSS.n394 2.77837
R8417 VSS.n4960 VSS.n809 2.77837
R8418 VSS.n5467 VSS.n57 2.77837
R8419 VSS.n2791 VSS.n2036 2.7666
R8420 VSS.n3098 VSS.n1993 2.7666
R8421 VSS.n3183 VSS.n1959 2.7666
R8422 VSS.n3979 VSS.n1911 2.7666
R8423 VSS.n4711 VSS.n1203 2.73369
R8424 VSS.n4715 VSS.n1194 2.73369
R8425 VSS.n4733 VSS.n4732 2.73369
R8426 VSS.n3972 VSS.n3971 2.73369
R8427 VSS.n4213 VSS.n4212 2.73369
R8428 VSS.n5254 VSS.n5253 2.73369
R8429 VSS.n5047 VSS.n5046 2.73369
R8430 VSS.n5009 VSS.n737 2.73369
R8431 VSS.n4421 VSS.n4420 2.73369
R8432 VSS.n2516 VSS.n2515 2.73369
R8433 VSS.n5420 VSS.n95 2.7239
R8434 VSS.n5207 VSS.n394 2.7239
R8435 VSS.n4954 VSS.n809 2.7239
R8436 VSS.n5468 VSS.n5467 2.7239
R8437 VSS.n2656 VSS.n2655 2.71236
R8438 VSS.n2629 VSS.n2586 2.71236
R8439 VSS.n2649 VSS.n2632 2.71236
R8440 VSS.n2648 VSS.n2633 2.71236
R8441 VSS.n2645 VSS.n2644 2.71236
R8442 VSS.n2639 VSS.n2634 2.71236
R8443 VSS.n2638 VSS.n2635 2.71236
R8444 VSS.n2752 VSS.n2042 2.71236
R8445 VSS.n2751 VSS.n2043 2.71236
R8446 VSS.n2759 VSS.n2036 2.71236
R8447 VSS.n2825 VSS.n2824 2.71236
R8448 VSS.n2798 VSS.n2031 2.71236
R8449 VSS.n2818 VSS.n2801 2.71236
R8450 VSS.n2817 VSS.n2802 2.71236
R8451 VSS.n2814 VSS.n2813 2.71236
R8452 VSS.n2808 VSS.n2803 2.71236
R8453 VSS.n2807 VSS.n2804 2.71236
R8454 VSS.n3058 VSS.n1999 2.71236
R8455 VSS.n3057 VSS.n2000 2.71236
R8456 VSS.n3065 VSS.n1993 2.71236
R8457 VSS.n3118 VSS.n1990 2.71236
R8458 VSS.n3119 VSS.n1989 2.71236
R8459 VSS.n3127 VSS.n3122 2.71236
R8460 VSS.n3126 VSS.n3123 2.71236
R8461 VSS.n3134 VSS.n1984 2.71236
R8462 VSS.n3135 VSS.n1983 2.71236
R8463 VSS.n3139 VSS.n3138 2.71236
R8464 VSS.n3144 VSS.n3141 2.71236
R8465 VSS.n3143 VSS.n3142 2.71236
R8466 VSS.n3151 VSS.n1959 2.71236
R8467 VSS.n3248 VSS.n3247 2.71236
R8468 VSS.n3190 VSS.n1955 2.71236
R8469 VSS.n3241 VSS.n3193 2.71236
R8470 VSS.n3240 VSS.n3194 2.71236
R8471 VSS.n3237 VSS.n3236 2.71236
R8472 VSS.n3199 VSS.n3195 2.71236
R8473 VSS.n3230 VSS.n3202 2.71236
R8474 VSS.n3229 VSS.n3227 2.71236
R8475 VSS.n3226 VSS.n3225 2.71236
R8476 VSS.n3979 VSS.n1913 2.71236
R8477 VSS.n4102 VSS.n4097 2.71236
R8478 VSS.n4101 VSS.n4098 2.71236
R8479 VSS.n4109 VSS.n1906 2.71236
R8480 VSS.n4110 VSS.n1905 2.71236
R8481 VSS.n4118 VSS.n4113 2.71236
R8482 VSS.n4117 VSS.n4114 2.71236
R8483 VSS.n4125 VSS.n1902 2.71236
R8484 VSS.n4128 VSS.n4127 2.71236
R8485 VSS.n4149 VSS.n4129 2.71236
R8486 VSS.n5375 VSS.n5374 2.64083
R8487 VSS.n8 VSS.n6 2.64083
R8488 VSS.n2299 VSS.n2298 2.61497
R8489 VSS.n2358 VSS.n2264 2.61497
R8490 VSS.n5421 VSS.n5419 2.61497
R8491 VSS.n5208 VSS.n5206 2.61497
R8492 VSS.n4955 VSS.n4953 2.61497
R8493 VSS.n5469 VSS.n62 2.61497
R8494 VSS.n5514 VSS.n5513 2.61497
R8495 VSS.n2370 VSS.n2264 2.61359
R8496 VSS.n2758 VSS.n2038 2.60389
R8497 VSS.n3064 VSS.n1995 2.60389
R8498 VSS.n3150 VSS.n1979 2.60389
R8499 VSS.n3221 VSS.n3220 2.60389
R8500 VSS.n4148 VSS.n1868 2.60389
R8501 VSS.n2683 VSS.n2682 2.59839
R8502 VSS.n4709 VSS.n1209 2.59839
R8503 VSS.n4767 VSS.n1129 2.59839
R8504 VSS.n4730 VSS.n1164 2.59839
R8505 VSS.n4073 VSS.n1833 2.59839
R8506 VSS.n5288 VSS.n267 2.59839
R8507 VSS.n5081 VSS.n302 2.59839
R8508 VSS.n5013 VSS.n730 2.59839
R8509 VSS.n4455 VSS.n742 2.59839
R8510 VSS.n4320 VSS.n1566 2.59839
R8511 VSS.n2306 VSS.n2277 2.58636
R8512 VSS.n2531 VSS.n2530 2.45707
R8513 VSS.n2551 VSS.n2251 2.45707
R8514 VSS.n2684 VSS.n2581 2.45707
R8515 VSS.n4211 VSS.n1853 2.45707
R8516 VSS.n1377 VSS.n1376 2.3255
R8517 VSS.n1375 VSS.n1371 2.3255
R8518 VSS.n5419 VSS.n5418 2.28816
R8519 VSS.n5206 VSS.n5205 2.28816
R8520 VSS.n4953 VSS.n4952 2.28816
R8521 VSS.n3645 VSS.n62 2.28816
R8522 VSS.n5514 VSS.n5512 2.28816
R8523 VSS.n2043 VSS.n2038 2.27847
R8524 VSS.n2000 VSS.n1995 2.27847
R8525 VSS.n3142 VSS.n1979 2.27847
R8526 VSS.n3225 VSS.n3221 2.27847
R8527 VSS.n4149 VSS.n4148 2.27847
R8528 VSS.n2656 VSS.n2585 2.16999
R8529 VSS.n2655 VSS.n2586 2.16999
R8530 VSS.n2632 VSS.n2629 2.16999
R8531 VSS.n2649 VSS.n2648 2.16999
R8532 VSS.n2645 VSS.n2633 2.16999
R8533 VSS.n2644 VSS.n2634 2.16999
R8534 VSS.n2639 VSS.n2638 2.16999
R8535 VSS.n2635 VSS.n2042 2.16999
R8536 VSS.n2752 VSS.n2751 2.16999
R8537 VSS.n2825 VSS.n2030 2.16999
R8538 VSS.n2824 VSS.n2031 2.16999
R8539 VSS.n2801 VSS.n2798 2.16999
R8540 VSS.n2818 VSS.n2817 2.16999
R8541 VSS.n2814 VSS.n2802 2.16999
R8542 VSS.n2813 VSS.n2803 2.16999
R8543 VSS.n2808 VSS.n2807 2.16999
R8544 VSS.n2804 VSS.n1999 2.16999
R8545 VSS.n3058 VSS.n3057 2.16999
R8546 VSS.n3110 VSS.n1990 2.16999
R8547 VSS.n3119 VSS.n3118 2.16999
R8548 VSS.n3122 VSS.n1989 2.16999
R8549 VSS.n3127 VSS.n3126 2.16999
R8550 VSS.n3123 VSS.n1984 2.16999
R8551 VSS.n3135 VSS.n3134 2.16999
R8552 VSS.n3138 VSS.n1983 2.16999
R8553 VSS.n3141 VSS.n3139 2.16999
R8554 VSS.n3144 VSS.n3143 2.16999
R8555 VSS.n3248 VSS.n1954 2.16999
R8556 VSS.n3247 VSS.n1955 2.16999
R8557 VSS.n3193 VSS.n3190 2.16999
R8558 VSS.n3241 VSS.n3240 2.16999
R8559 VSS.n3237 VSS.n3194 2.16999
R8560 VSS.n3236 VSS.n3195 2.16999
R8561 VSS.n3202 VSS.n3199 2.16999
R8562 VSS.n3230 VSS.n3229 2.16999
R8563 VSS.n3227 VSS.n3226 2.16999
R8564 VSS.n4097 VSS.n1910 2.16999
R8565 VSS.n4102 VSS.n4101 2.16999
R8566 VSS.n4098 VSS.n1906 2.16999
R8567 VSS.n4110 VSS.n4109 2.16999
R8568 VSS.n4113 VSS.n1905 2.16999
R8569 VSS.n4118 VSS.n4117 2.16999
R8570 VSS.n4114 VSS.n1902 2.16999
R8571 VSS.n4127 VSS.n4125 2.16999
R8572 VSS.n4129 VSS.n4128 2.16999
R8573 VSS.n1224 VSS.n1223 2.12075
R8574 VSS.n1275 VSS.n1056 2.12075
R8575 VSS.n4010 VSS.n1780 2.12075
R8576 VSS.n3924 VSS.n3867 2.12075
R8577 VSS.n5368 VSS.n123 2.07029
R8578 VSS.n5159 VSS.n5158 2.07029
R8579 VSS.n4906 VSS.n4905 2.07029
R8580 VSS.n3623 VSS.n3622 2.07029
R8581 VSS.n5479 VSS.n5478 2.07029
R8582 VSS.n2585 VSS.n2584 2.06152
R8583 VSS.n2030 VSS.n2029 2.06152
R8584 VSS.n3111 VSS.n3110 2.06152
R8585 VSS.n1954 VSS.n1953 2.06152
R8586 VSS.n4081 VSS.n1910 2.06152
R8587 VSS.n4631 VSS.n1397 1.89388
R8588 VSS.n4635 VSS.n1394 1.86266
R8589 VSS.n4637 VSS.n4636 1.8605
R8590 VSS.n4634 VSS.n4633 1.8605
R8591 VSS.n4686 VSS.n1224 1.8459
R8592 VSS.n1340 VSS.n1056 1.8459
R8593 VSS.n4014 VSS.n1780 1.8459
R8594 VSS.n3924 VSS.n3923 1.8459
R8595 VSS.n4190 VSS.n1357 1.80664
R8596 VSS.n4595 VSS.n24 1.77399
R8597 VSS.n2572 VSS.n2239 1.76337
R8598 VSS.n4644 VSS.n1387 1.76337
R8599 VSS.n5536 VSS.n22 1.61978
R8600 VSS.n1899 VSS.n1898 1.52394
R8601 VSS VSS.n1877 1.46383
R8602 VSS.n4584 VSS.n1387 1.45679
R8603 VSS.n2298 VSS.n168 1.41667
R8604 VSS.n1880 VSS 1.41317
R8605 VSS.n2682 VSS.n2675 1.40769
R8606 VSS.n2848 VSS.n1209 1.40769
R8607 VSS.n4768 VSS.n4767 1.40769
R8608 VSS.n3271 VSS.n1164 1.40769
R8609 VSS.n4273 VSS.n1833 1.40769
R8610 VSS.n5289 VSS.n5288 1.40769
R8611 VSS.n5082 VSS.n5081 1.40769
R8612 VSS.n4829 VSS.n730 1.40769
R8613 VSS.n4456 VSS.n4455 1.40769
R8614 VSS.n4321 VSS.n4320 1.40769
R8615 VSS.n2358 VSS.n2357 1.38944
R8616 VSS.n4710 VSS.n4709 1.38063
R8617 VSS.n1196 VSS.n1129 1.38063
R8618 VSS.n4731 VSS.n4730 1.38063
R8619 VSS.n4073 VSS.n3998 1.38063
R8620 VSS.n302 VSS.n299 1.38063
R8621 VSS.n5013 VSS.n727 1.38063
R8622 VSS.n742 VSS.n740 1.38063
R8623 VSS.n1566 VSS.n1563 1.38063
R8624 VSS.n4711 VSS.n4710 1.35357
R8625 VSS.n4715 VSS.n1196 1.35357
R8626 VSS.n4732 VSS.n4731 1.35357
R8627 VSS.n3998 VSS.n3972 1.35357
R8628 VSS.n5253 VSS.n299 1.35357
R8629 VSS.n5046 VSS.n727 1.35357
R8630 VSS.n5009 VSS.n740 1.35357
R8631 VSS.n4420 VSS.n1563 1.35357
R8632 VSS.n2121 VSS.n1203 1.29944
R8633 VSS.n2900 VSS.n1194 1.29944
R8634 VSS.n4733 VSS.n1153 1.29944
R8635 VSS.n3971 VSS.n1922 1.29944
R8636 VSS.n4213 VSS.n1849 1.29944
R8637 VSS.n5254 VSS.n291 1.29944
R8638 VSS.n5047 VSS.n719 1.29944
R8639 VSS.n3811 VSS.n737 1.29944
R8640 VSS.n4421 VSS.n1556 1.29944
R8641 VSS.n2515 VSS.n2409 1.29944
R8642 VSS.n5467 VSS.n5466 1.29343
R8643 VSS.n394 VSS.n393 1.29343
R8644 VSS.n809 VSS.n808 1.29343
R8645 VSS.n153 VSS.n95 1.29343
R8646 VSS.n4633 VSS 1.28778
R8647 VSS.n1234 VSS.n299 1.22878
R8648 VSS.n1314 VSS.n727 1.22878
R8649 VSS.n4044 VSS.n1563 1.22878
R8650 VSS.n3881 VSS.n740 1.22878
R8651 VSS.n3998 VSS.n3997 1.22878
R8652 VSS.n3093 VSS.n1196 1.22878
R8653 VSS.n4731 VSS.n1162 1.22878
R8654 VSS.n4710 VSS.n1207 1.22878
R8655 VSS VSS.n0 1.16168
R8656 VSS.n595 VSS.n594 1.14433
R8657 VSS.n638 VSS.n637 1.14433
R8658 VSS.n962 VSS.n961 1.14433
R8659 VSS.n4583 VSS.n1407 1.14433
R8660 VSS.n5532 VSS.n5531 1.14433
R8661 VSS.n4501 VSS.n1453 1.14433
R8662 VSS.n1650 VSS.n1649 1.14433
R8663 VSS.n3684 VSS.n3449 1.14433
R8664 VSS.n3736 VSS.n3735 1.14433
R8665 VSS.n941 VSS.n940 1.14433
R8666 VSS.n2986 VSS.n2985 1.13948
R8667 VSS.n2207 VSS.n2206 1.13948
R8668 VSS.n3383 VSS.n3382 1.13948
R8669 VSS.n3866 VSS.n3865 1.13948
R8670 VSS.n2490 VSS.n2489 1.13948
R8671 VSS.n2160 VSS.n2121 1.13708
R8672 VSS.n2939 VSS.n2900 1.13708
R8673 VSS.n4737 VSS.n1153 1.13708
R8674 VSS.n3967 VSS.n1922 1.13708
R8675 VSS.n4217 VSS.n1849 1.13708
R8676 VSS.n5258 VSS.n291 1.13708
R8677 VSS.n5051 VSS.n719 1.13708
R8678 VSS.n3811 VSS.n3810 1.13708
R8679 VSS.n4425 VSS.n1556 1.13708
R8680 VSS.n2511 VSS.n2409 1.13708
R8681 VSS.n5349 VSS.n169 1.08986
R8682 VSS.n173 VSS.n170 1.08986
R8683 VSS.n5344 VSS.n176 1.08986
R8684 VSS.n5334 VSS.n178 1.08986
R8685 VSS.n5338 VSS.n5337 1.08986
R8686 VSS.n580 VSS.n579 1.08986
R8687 VSS.n586 VSS.n584 1.08986
R8688 VSS.n589 VSS.n588 1.08986
R8689 VSS.n5329 VSS.n202 1.08986
R8690 VSS.n206 VSS.n203 1.08986
R8691 VSS.n5324 VSS.n207 1.08986
R8692 VSS.n215 VSS.n210 1.08986
R8693 VSS.n5318 VSS.n5317 1.08986
R8694 VSS.n624 VSS.n218 1.08986
R8695 VSS.n627 VSS.n622 1.08986
R8696 VSS.n632 VSS.n631 1.08986
R8697 VSS.n5139 VSS.n423 1.08986
R8698 VSS.n427 VSS.n424 1.08986
R8699 VSS.n5134 VSS.n430 1.08986
R8700 VSS.n5130 VSS.n5129 1.08986
R8701 VSS.n5126 VSS.n438 1.08986
R8702 VSS.n862 VSS.n851 1.08986
R8703 VSS.n868 VSS.n867 1.08986
R8704 VSS.n873 VSS.n872 1.08986
R8705 VSS.n4398 VSS.n4397 1.08986
R8706 VSS.n1693 VSS.n1690 1.08986
R8707 VSS.n4375 VSS.n1696 1.08986
R8708 VSS.n4365 VSS.n1699 1.08986
R8709 VSS.n4369 VSS.n4368 1.08986
R8710 VSS.n1722 VSS.n1713 1.08986
R8711 VSS.n1728 VSS.n1727 1.08986
R8712 VSS.n1736 VSS.n1735 1.08986
R8713 VSS.n4505 VSS.n1444 1.08986
R8714 VSS.n4576 VSS.n1445 1.08986
R8715 VSS.n4572 VSS.n4571 1.08986
R8716 VSS.n4567 VSS.n4529 1.08986
R8717 VSS.n4563 VSS.n4530 1.08986
R8718 VSS.n4557 VSS.n4556 1.08986
R8719 VSS.n4552 VSS.n4543 1.08986
R8720 VSS.n4548 VSS.n4544 1.08986
R8721 VSS.n3486 VSS.n3479 1.08986
R8722 VSS.n3674 VSS.n3673 1.08986
R8723 VSS.n3523 VSS.n3522 1.08986
R8724 VSS.n3527 VSS.n3521 1.08986
R8725 VSS.n3532 VSS.n3518 1.08986
R8726 VSS.n3536 VSS.n3517 1.08986
R8727 VSS.n3549 VSS.n3548 1.08986
R8728 VSS.n3545 VSS.n3539 1.08986
R8729 VSS.n4494 VSS.n1475 1.08986
R8730 VSS.n1479 VSS.n1476 1.08986
R8731 VSS.n4489 VSS.n1481 1.08986
R8732 VSS.n4485 VSS.n4484 1.08986
R8733 VSS.n4481 VSS.n1489 1.08986
R8734 VSS.n1635 VSS.n1634 1.08986
R8735 VSS.n1640 VSS.n1639 1.08986
R8736 VSS.n1644 VSS.n1643 1.08986
R8737 VSS.n4886 VSS.n838 1.08986
R8738 VSS.n842 VSS.n839 1.08986
R8739 VSS.n4881 VSS.n845 1.08986
R8740 VSS.n4877 VSS.n4876 1.08986
R8741 VSS.n4873 VSS.n976 1.08986
R8742 VSS.n3464 VSS.n3454 1.08986
R8743 VSS.n3468 VSS.n3453 1.08986
R8744 VSS.n3473 VSS.n3450 1.08986
R8745 VSS.n4867 VSS.n996 1.08986
R8746 VSS.n1000 VSS.n997 1.08986
R8747 VSS.n4862 VSS.n1002 1.08986
R8748 VSS.n4858 VSS.n4857 1.08986
R8749 VSS.n4854 VSS.n1010 1.08986
R8750 VSS.n3721 VSS.n3720 1.08986
R8751 VSS.n3726 VSS.n3725 1.08986
R8752 VSS.n3730 VSS.n3729 1.08986
R8753 VSS.n5120 VSS.n458 1.08986
R8754 VSS.n462 VSS.n459 1.08986
R8755 VSS.n5115 VSS.n464 1.08986
R8756 VSS.n5111 VSS.n5110 1.08986
R8757 VSS.n5107 VSS.n469 1.08986
R8758 VSS.n926 VSS.n925 1.08986
R8759 VSS.n931 VSS.n930 1.08986
R8760 VSS.n935 VSS.n934 1.08986
R8761 VSS.n3018 VSS.n2856 1.08525
R8762 VSS.n3022 VSS.n3016 1.08525
R8763 VSS.n3013 VSS.n2858 1.08525
R8764 VSS.n2864 VSS.n2862 1.08525
R8765 VSS.n3007 VSS.n2867 1.08525
R8766 VSS.n2999 VSS.n2869 1.08525
R8767 VSS.n2876 VSS.n2873 1.08525
R8768 VSS.n2990 VSS.n2877 1.08525
R8769 VSS.n2712 VSS.n2079 1.08525
R8770 VSS.n2716 VSS.n2238 1.08525
R8771 VSS.n2235 VSS.n2081 1.08525
R8772 VSS.n2087 VSS.n2085 1.08525
R8773 VSS.n2229 VSS.n2090 1.08525
R8774 VSS.n2221 VSS.n2092 1.08525
R8775 VSS.n2099 VSS.n2096 1.08525
R8776 VSS.n2212 VSS.n2209 1.08525
R8777 VSS.n3926 VSS.n3279 1.08525
R8778 VSS.n3930 VSS.n3413 1.08525
R8779 VSS.n3410 VSS.n3281 1.08525
R8780 VSS.n3287 VSS.n3285 1.08525
R8781 VSS.n3404 VSS.n3290 1.08525
R8782 VSS.n3396 VSS.n3292 1.08525
R8783 VSS.n3299 VSS.n3296 1.08525
R8784 VSS.n3387 VSS.n3300 1.08525
R8785 VSS.n4791 VSS.n1058 1.08525
R8786 VSS.n4787 VSS.n4786 1.08525
R8787 VSS.n4783 VSS.n1064 1.08525
R8788 VSS.n3839 VSS.n1065 1.08525
R8789 VSS.n3843 VSS.n3842 1.08525
R8790 VSS.n3852 VSS.n3851 1.08525
R8791 VSS.n3858 VSS.n3856 1.08525
R8792 VSS.n3861 VSS.n3860 1.08525
R8793 VSS.n4295 VSS.n1782 1.08525
R8794 VSS.n4291 VSS.n4290 1.08525
R8795 VSS.n4287 VSS.n1785 1.08525
R8796 VSS.n2461 VSS.n1789 1.08525
R8797 VSS.n2465 VSS.n2464 1.08525
R8798 VSS.n2474 VSS.n2473 1.08525
R8799 VSS.n2481 VSS.n2478 1.08525
R8800 VSS.n2484 VSS.n2453 1.08525
R8801 VSS.n2678 VSS.n2064 1.08295
R8802 VSS.n2746 VSS.n2065 1.08295
R8803 VSS.n2742 VSS.n2741 1.08295
R8804 VSS.n2135 VSS.n2134 1.08295
R8805 VSS.n2140 VSS.n2127 1.08295
R8806 VSS.n2151 VSS.n2150 1.08295
R8807 VSS.n2165 VSS.n2124 1.08295
R8808 VSS.n2125 VSS.n2122 1.08295
R8809 VSS.n2847 VSS.n2021 1.08295
R8810 VSS.n3052 VSS.n2022 1.08295
R8811 VSS.n3048 VSS.n3047 1.08295
R8812 VSS.n2914 VSS.n2913 1.08295
R8813 VSS.n2919 VSS.n2906 1.08295
R8814 VSS.n2930 VSS.n2929 1.08295
R8815 VSS.n2944 VSS.n2903 1.08295
R8816 VSS.n2904 VSS.n2901 1.08295
R8817 VSS.n4778 VSS.n1088 1.08295
R8818 VSS.n1092 VSS.n1089 1.08295
R8819 VSS.n4759 VSS.n4758 1.08295
R8820 VSS.n4755 VSS.n1135 1.08295
R8821 VSS.n1137 VSS.n1136 1.08295
R8822 VSS.n4746 VSS.n4745 1.08295
R8823 VSS.n4742 VSS.n1150 1.08295
R8824 VSS.n1152 VSS.n1151 1.08295
R8825 VSS.n3270 VSS.n1945 1.08295
R8826 VSS.n3960 VSS.n1946 1.08295
R8827 VSS.n3956 VSS.n3955 1.08295
R8828 VSS.n3317 VSS.n3316 1.08295
R8829 VSS.n3322 VSS.n3309 1.08295
R8830 VSS.n3333 VSS.n3332 1.08295
R8831 VSS.n3341 VSS.n3307 1.08295
R8832 VSS.n3339 VSS.n1924 1.08295
R8833 VSS.n4256 VSS.n1835 1.08295
R8834 VSS.n4279 VSS.n1810 1.08295
R8835 VSS.n1838 VSS.n1811 1.08295
R8836 VSS.n4242 VSS.n1840 1.08295
R8837 VSS.n4246 VSS.n4245 1.08295
R8838 VSS.n4234 VSS.n4233 1.08295
R8839 VSS.n4226 VSS.n1846 1.08295
R8840 VSS.n4222 VSS.n4221 1.08295
R8841 VSS.n5309 VSS.n241 1.08295
R8842 VSS.n245 VSS.n242 1.08295
R8843 VSS.n5280 VSS.n5279 1.08295
R8844 VSS.n5276 VSS.n273 1.08295
R8845 VSS.n275 VSS.n274 1.08295
R8846 VSS.n5267 VSS.n5266 1.08295
R8847 VSS.n5263 VSS.n288 1.08295
R8848 VSS.n290 VSS.n289 1.08295
R8849 VSS.n5102 VSS.n490 1.08295
R8850 VSS.n494 VSS.n491 1.08295
R8851 VSS.n5073 VSS.n5072 1.08295
R8852 VSS.n5069 VSS.n701 1.08295
R8853 VSS.n703 VSS.n702 1.08295
R8854 VSS.n5060 VSS.n5059 1.08295
R8855 VSS.n5056 VSS.n716 1.08295
R8856 VSS.n718 VSS.n717 1.08295
R8857 VSS.n4849 VSS.n1031 1.08295
R8858 VSS.n1035 VSS.n1032 1.08295
R8859 VSS.n3779 VSS.n3777 1.08295
R8860 VSS.n3782 VSS.n3759 1.08295
R8861 VSS.n3787 VSS.n3758 1.08295
R8862 VSS.n3795 VSS.n3757 1.08295
R8863 VSS.n3798 VSS.n3756 1.08295
R8864 VSS.n3805 VSS.n3804 1.08295
R8865 VSS.n4476 VSS.n1510 1.08295
R8866 VSS.n1514 VSS.n1511 1.08295
R8867 VSS.n4447 VSS.n4446 1.08295
R8868 VSS.n4443 VSS.n1538 1.08295
R8869 VSS.n1540 VSS.n1539 1.08295
R8870 VSS.n4434 VSS.n4433 1.08295
R8871 VSS.n4430 VSS.n1553 1.08295
R8872 VSS.n1555 VSS.n1554 1.08295
R8873 VSS.n4359 VSS.n1751 1.08295
R8874 VSS.n1755 VSS.n1752 1.08295
R8875 VSS.n4354 VSS.n1757 1.08295
R8876 VSS.n4344 VSS.n1759 1.08295
R8877 VSS.n4348 VSS.n4347 1.08295
R8878 VSS.n2426 VSS.n2413 1.08295
R8879 VSS.n2431 VSS.n2412 1.08295
R8880 VSS.n2434 VSS.n2411 1.08295
R8881 VSS.n4631 VSS 1.07635
R8882 VSS.n576 VSS 1.06263
R8883 VSS.n5314 VSS 1.06263
R8884 VSS.n859 VSS 1.06263
R8885 VSS.n1719 VSS 1.06263
R8886 VSS.n4540 VSS 1.06263
R8887 VSS.n3560 VSS 1.06263
R8888 VSS.n1631 VSS 1.06263
R8889 VSS.n3462 VSS 1.06263
R8890 VSS.n3717 VSS 1.06263
R8891 VSS.n922 VSS 1.06263
R8892 VSS VSS.n3002 1.05813
R8893 VSS VSS.n2224 1.05813
R8894 VSS VSS.n3399 1.05813
R8895 VSS.n3848 VSS 1.05813
R8896 VSS.n2470 VSS 1.05813
R8897 VSS.n2145 VSS 1.05589
R8898 VSS.n2924 VSS 1.05589
R8899 VSS.n1145 VSS 1.05589
R8900 VSS.n3327 VSS 1.05589
R8901 VSS.n4230 VSS 1.05589
R8902 VSS.n283 VSS 1.05589
R8903 VSS.n711 VSS 1.05589
R8904 VSS.n3790 VSS 1.05589
R8905 VSS.n1548 VSS 1.05589
R8906 VSS.n2423 VSS 1.05589
R8907 VSS.n169 VSS.n168 1.03539
R8908 VSS.n2356 VSS.n202 1.03539
R8909 VSS.n423 VSS.n422 1.03539
R8910 VSS.n4398 VSS.n1689 1.03539
R8911 VSS.n4506 VSS.n4505 1.03539
R8912 VSS.n3604 VSS.n3479 1.03539
R8913 VSS.n3586 VSS.n1475 1.03539
R8914 VSS.n838 VSS.n837 1.03539
R8915 VSS.n4811 VSS.n996 1.03539
R8916 VSS.n680 VSS.n458 1.03539
R8917 VSS.n3018 VSS.n3017 1.03101
R8918 VSS.n2712 VSS.n2711 1.03101
R8919 VSS.n3926 VSS.n3925 1.03101
R8920 VSS.n4792 VSS.n4791 1.03101
R8921 VSS.n4296 VSS.n4295 1.03101
R8922 VSS.n2678 VSS.n2675 1.02883
R8923 VSS.n2848 VSS.n2847 1.02883
R8924 VSS.n4768 VSS.n1088 1.02883
R8925 VSS.n3271 VSS.n3270 1.02883
R8926 VSS.n4273 VSS.n4256 1.02883
R8927 VSS.n5289 VSS.n241 1.02883
R8928 VSS.n5082 VSS.n490 1.02883
R8929 VSS.n4829 VSS.n1031 1.02883
R8930 VSS.n4456 VSS.n1510 1.02883
R8931 VSS.n4321 VSS.n1751 1.02883
R8932 VSS.n595 VSS.n83 0.980926
R8933 VSS.n679 VSS.n638 0.980926
R8934 VSS.n422 VSS.n83 0.980926
R8935 VSS.n961 VSS.n847 0.980926
R8936 VSS.n1689 VSS.n1651 0.980926
R8937 VSS.n4584 VSS.n4583 0.980926
R8938 VSS.n4506 VSS.n4502 0.980926
R8939 VSS.n5531 VSS.n22 0.980926
R8940 VSS.n3604 VSS.n3478 0.980926
R8941 VSS.n4502 VSS.n4501 0.980926
R8942 VSS.n3586 VSS.n761 0.980926
R8943 VSS.n1651 VSS.n1650 0.980926
R8944 VSS.n847 VSS.n837 0.980926
R8945 VSS.n3478 VSS.n3449 0.980926
R8946 VSS.n4811 VSS.n332 0.980926
R8947 VSS.n3736 VSS.n761 0.980926
R8948 VSS.n680 VSS.n679 0.980926
R8949 VSS.n941 VSS.n332 0.980926
R8950 VSS.n3017 VSS.n1224 0.976771
R8951 VSS.n2985 VSS.n1056 0.976771
R8952 VSS.n2711 VSS.n2710 0.976771
R8953 VSS.n2206 VSS.n1224 0.976771
R8954 VSS.n3925 VSS.n3924 0.976771
R8955 VSS.n3382 VSS.n1780 0.976771
R8956 VSS.n4792 VSS.n1056 0.976771
R8957 VSS.n3924 VSS.n3866 0.976771
R8958 VSS.n4296 VSS.n1780 0.976771
R8959 VSS.n2490 VSS.n1360 0.976771
R8960 VSS.n5349 VSS.n5348 0.926457
R8961 VSS.n5345 VSS.n173 0.926457
R8962 VSS.n182 VSS.n176 0.926457
R8963 VSS.n5334 VSS.n180 0.926457
R8964 VSS.n5337 VSS.n5333 0.926457
R8965 VSS.n576 VSS.n573 0.926457
R8966 VSS.n579 VSS.n571 0.926457
R8967 VSS.n587 VSS.n586 0.926457
R8968 VSS.n588 VSS.n568 0.926457
R8969 VSS.n5329 VSS.n5328 0.926457
R8970 VSS.n5325 VSS.n206 0.926457
R8971 VSS.n223 VSS.n207 0.926457
R8972 VSS.n216 VSS.n215 0.926457
R8973 VSS.n5317 VSS.n217 0.926457
R8974 VSS.n5314 VSS.n5313 0.926457
R8975 VSS.n624 VSS.n623 0.926457
R8976 VSS.n628 VSS.n627 0.926457
R8977 VSS.n631 VSS.n614 0.926457
R8978 VSS.n5139 VSS.n5138 0.926457
R8979 VSS.n5135 VSS.n427 0.926457
R8980 VSS.n436 VSS.n430 0.926457
R8981 VSS.n5129 VSS.n437 0.926457
R8982 VSS.n5126 VSS.n5125 0.926457
R8983 VSS.n859 VSS.n858 0.926457
R8984 VSS.n865 VSS.n862 0.926457
R8985 VSS.n867 VSS.n849 0.926457
R8986 VSS.n874 VSS.n873 0.926457
R8987 VSS.n4397 VSS.n4379 0.926457
R8988 VSS.n4376 VSS.n1693 0.926457
R8989 VSS.n1703 VSS.n1696 0.926457
R8990 VSS.n4365 VSS.n1701 0.926457
R8991 VSS.n4368 VSS.n4364 0.926457
R8992 VSS.n1719 VSS.n1718 0.926457
R8993 VSS.n1725 VSS.n1722 0.926457
R8994 VSS.n1727 VSS.n1711 0.926457
R8995 VSS.n1737 VSS.n1736 0.926457
R8996 VSS.n4577 VSS.n1444 0.926457
R8997 VSS.n1448 VSS.n1445 0.926457
R8998 VSS.n4571 VSS.n1449 0.926457
R8999 VSS.n4567 VSS.n4566 0.926457
R9000 VSS.n4535 VSS.n4530 0.926457
R9001 VSS.n4540 VSS.n4538 0.926457
R9002 VSS.n4556 VSS.n4539 0.926457
R9003 VSS.n4552 VSS.n4551 0.926457
R9004 VSS.n4544 VSS.n27 0.926457
R9005 VSS.n3486 VSS.n3481 0.926457
R9006 VSS.n3673 VSS.n3484 0.926457
R9007 VSS.n3528 VSS.n3522 0.926457
R9008 VSS.n3531 VSS.n3521 0.926457
R9009 VSS.n3556 VSS.n3518 0.926457
R9010 VSS.n3560 VSS.n3559 0.926457
R9011 VSS.n3538 VSS.n3536 0.926457
R9012 VSS.n3548 VSS.n3546 0.926457
R9013 VSS.n3539 VSS.n1456 0.926457
R9014 VSS.n4494 VSS.n4493 0.926457
R9015 VSS.n4490 VSS.n1479 0.926457
R9016 VSS.n1487 VSS.n1481 0.926457
R9017 VSS.n4484 VSS.n1488 0.926457
R9018 VSS.n4481 VSS.n4480 0.926457
R9019 VSS.n1631 VSS.n1626 0.926457
R9020 VSS.n1634 VSS.n1624 0.926457
R9021 VSS.n1640 VSS.n1622 0.926457
R9022 VSS.n1643 VSS.n1620 0.926457
R9023 VSS.n4886 VSS.n4885 0.926457
R9024 VSS.n4882 VSS.n842 0.926457
R9025 VSS.n974 VSS.n845 0.926457
R9026 VSS.n4876 VSS.n975 0.926457
R9027 VSS.n4873 VSS.n4872 0.926457
R9028 VSS.n3463 VSS.n3462 0.926457
R9029 VSS.n3469 VSS.n3454 0.926457
R9030 VSS.n3472 VSS.n3453 0.926457
R9031 VSS.n3685 VSS.n3450 0.926457
R9032 VSS.n4867 VSS.n4866 0.926457
R9033 VSS.n4863 VSS.n1000 0.926457
R9034 VSS.n1008 VSS.n1002 0.926457
R9035 VSS.n4857 VSS.n1009 0.926457
R9036 VSS.n4854 VSS.n4853 0.926457
R9037 VSS.n3717 VSS.n3712 0.926457
R9038 VSS.n3720 VSS.n3710 0.926457
R9039 VSS.n3726 VSS.n3708 0.926457
R9040 VSS.n3729 VSS.n3706 0.926457
R9041 VSS.n5120 VSS.n5119 0.926457
R9042 VSS.n5116 VSS.n462 0.926457
R9043 VSS.n467 VSS.n464 0.926457
R9044 VSS.n5110 VSS.n468 0.926457
R9045 VSS.n5107 VSS.n5106 0.926457
R9046 VSS.n922 VSS.n917 0.926457
R9047 VSS.n925 VSS.n915 0.926457
R9048 VSS.n931 VSS.n913 0.926457
R9049 VSS.n934 VSS.n911 0.926457
R9050 VSS.n3023 VSS.n2856 0.922534
R9051 VSS.n3016 VSS.n2857 0.922534
R9052 VSS.n3013 VSS.n3012 0.922534
R9053 VSS.n3008 VSS.n2864 0.922534
R9054 VSS.n2993 VSS.n2867 0.922534
R9055 VSS.n3002 VSS.n2868 0.922534
R9056 VSS.n2999 VSS.n2998 0.922534
R9057 VSS.n2991 VSS.n2876 0.922534
R9058 VSS.n2878 VSS.n2877 0.922534
R9059 VSS.n2717 VSS.n2079 0.922534
R9060 VSS.n2238 VSS.n2080 0.922534
R9061 VSS.n2235 VSS.n2234 0.922534
R9062 VSS.n2230 VSS.n2087 0.922534
R9063 VSS.n2215 VSS.n2090 0.922534
R9064 VSS.n2224 VSS.n2091 0.922534
R9065 VSS.n2221 VSS.n2220 0.922534
R9066 VSS.n2213 VSS.n2099 0.922534
R9067 VSS.n2209 VSS.n2208 0.922534
R9068 VSS.n3931 VSS.n3279 0.922534
R9069 VSS.n3413 VSS.n3280 0.922534
R9070 VSS.n3410 VSS.n3409 0.922534
R9071 VSS.n3405 VSS.n3287 0.922534
R9072 VSS.n3390 VSS.n3290 0.922534
R9073 VSS.n3399 VSS.n3291 0.922534
R9074 VSS.n3396 VSS.n3395 0.922534
R9075 VSS.n3388 VSS.n3299 0.922534
R9076 VSS.n3301 VSS.n3300 0.922534
R9077 VSS.n1062 VSS.n1058 0.922534
R9078 VSS.n4786 VSS.n1063 0.922534
R9079 VSS.n4783 VSS.n4782 0.922534
R9080 VSS.n3839 VSS.n3835 0.922534
R9081 VSS.n3842 VSS.n3838 0.922534
R9082 VSS.n3848 VSS.n3834 0.922534
R9083 VSS.n3851 VSS.n3833 0.922534
R9084 VSS.n3859 VSS.n3858 0.922534
R9085 VSS.n3860 VSS.n3831 0.922534
R9086 VSS.n1783 VSS.n1782 0.922534
R9087 VSS.n4290 VSS.n1784 0.922534
R9088 VSS.n4287 VSS.n4286 0.922534
R9089 VSS.n2461 VSS.n2458 0.922534
R9090 VSS.n2464 VSS.n2460 0.922534
R9091 VSS.n2470 VSS.n2457 0.922534
R9092 VSS.n2473 VSS.n2454 0.922534
R9093 VSS.n2485 VSS.n2481 0.922534
R9094 VSS.n2488 VSS.n2453 0.922534
R9095 VSS.n2747 VSS.n2064 0.920585
R9096 VSS.n2068 VSS.n2065 0.920585
R9097 VSS.n2741 VSS.n2070 0.920585
R9098 VSS.n2136 VSS.n2135 0.920585
R9099 VSS.n2140 VSS.n2139 0.920585
R9100 VSS.n2146 VSS.n2145 0.920585
R9101 VSS.n2150 VSS.n2149 0.920585
R9102 VSS.n2165 VSS.n2164 0.920585
R9103 VSS.n2161 VSS.n2122 0.920585
R9104 VSS.n3053 VSS.n2021 0.920585
R9105 VSS.n2025 VSS.n2022 0.920585
R9106 VSS.n3047 VSS.n2027 0.920585
R9107 VSS.n2915 VSS.n2914 0.920585
R9108 VSS.n2919 VSS.n2918 0.920585
R9109 VSS.n2925 VSS.n2924 0.920585
R9110 VSS.n2929 VSS.n2928 0.920585
R9111 VSS.n2944 VSS.n2943 0.920585
R9112 VSS.n2940 VSS.n2901 0.920585
R9113 VSS.n4778 VSS.n4777 0.920585
R9114 VSS.n1093 VSS.n1092 0.920585
R9115 VSS.n4758 VSS.n1134 0.920585
R9116 VSS.n4755 VSS.n4754 0.920585
R9117 VSS.n4751 VSS.n1137 0.920585
R9118 VSS.n1146 VSS.n1145 0.920585
R9119 VSS.n4745 VSS.n1149 0.920585
R9120 VSS.n4742 VSS.n4741 0.920585
R9121 VSS.n4738 VSS.n1152 0.920585
R9122 VSS.n3961 VSS.n1945 0.920585
R9123 VSS.n1949 VSS.n1946 0.920585
R9124 VSS.n3955 VSS.n1951 0.920585
R9125 VSS.n3318 VSS.n3317 0.920585
R9126 VSS.n3322 VSS.n3321 0.920585
R9127 VSS.n3328 VSS.n3327 0.920585
R9128 VSS.n3332 VSS.n3331 0.920585
R9129 VSS.n3341 VSS.n3340 0.920585
R9130 VSS.n3966 VSS.n1924 0.920585
R9131 VSS.n1835 VSS.n1834 0.920585
R9132 VSS.n4279 VSS.n4278 0.920585
R9133 VSS.n1839 VSS.n1838 0.920585
R9134 VSS.n4242 VSS.n1842 0.920585
R9135 VSS.n4245 VSS.n4241 0.920585
R9136 VSS.n4230 VSS.n1844 0.920585
R9137 VSS.n4233 VSS.n4229 0.920585
R9138 VSS.n1848 VSS.n1846 0.920585
R9139 VSS.n4221 VSS.n4220 0.920585
R9140 VSS.n5309 VSS.n5308 0.920585
R9141 VSS.n246 VSS.n245 0.920585
R9142 VSS.n5279 VSS.n272 0.920585
R9143 VSS.n5276 VSS.n5275 0.920585
R9144 VSS.n5272 VSS.n275 0.920585
R9145 VSS.n284 VSS.n283 0.920585
R9146 VSS.n5266 VSS.n287 0.920585
R9147 VSS.n5263 VSS.n5262 0.920585
R9148 VSS.n5259 VSS.n290 0.920585
R9149 VSS.n5102 VSS.n5101 0.920585
R9150 VSS.n495 VSS.n494 0.920585
R9151 VSS.n5072 VSS.n700 0.920585
R9152 VSS.n5069 VSS.n5068 0.920585
R9153 VSS.n5065 VSS.n703 0.920585
R9154 VSS.n712 VSS.n711 0.920585
R9155 VSS.n5059 VSS.n715 0.920585
R9156 VSS.n5056 VSS.n5055 0.920585
R9157 VSS.n5052 VSS.n718 0.920585
R9158 VSS.n4849 VSS.n4848 0.920585
R9159 VSS.n1036 VSS.n1035 0.920585
R9160 VSS.n3779 VSS.n3778 0.920585
R9161 VSS.n3783 VSS.n3782 0.920585
R9162 VSS.n3787 VSS.n3786 0.920585
R9163 VSS.n3791 VSS.n3790 0.920585
R9164 VSS.n3795 VSS.n3794 0.920585
R9165 VSS.n3801 VSS.n3798 0.920585
R9166 VSS.n3804 VSS.n3754 0.920585
R9167 VSS.n4476 VSS.n4475 0.920585
R9168 VSS.n1515 VSS.n1514 0.920585
R9169 VSS.n4446 VSS.n1537 0.920585
R9170 VSS.n4443 VSS.n4442 0.920585
R9171 VSS.n4439 VSS.n1540 0.920585
R9172 VSS.n1549 VSS.n1548 0.920585
R9173 VSS.n4433 VSS.n1552 0.920585
R9174 VSS.n4430 VSS.n4429 0.920585
R9175 VSS.n4426 VSS.n1555 0.920585
R9176 VSS.n4359 VSS.n4358 0.920585
R9177 VSS.n4355 VSS.n1755 0.920585
R9178 VSS.n4338 VSS.n1757 0.920585
R9179 VSS.n4344 VSS.n1761 0.920585
R9180 VSS.n4347 VSS.n4343 0.920585
R9181 VSS.n2423 VSS.n2422 0.920585
R9182 VSS.n2427 VSS.n2426 0.920585
R9183 VSS.n2431 VSS.n2430 0.920585
R9184 VSS.n2510 VSS.n2434 0.920585
R9185 VSS.n4403 VSS.n4402 0.903568
R9186 VSS.n1451 VSS.n74 0.903568
R9187 VSS.n4992 VSS.n4991 0.903568
R9188 VSS.n5232 VSS.n5231 0.903568
R9189 VSS.n846 VSS.n359 0.903568
R9190 VSS.n3477 VSS.n3476 0.903568
R9191 VSS.n5434 VSS.n5433 0.903568
R9192 VSS.n5236 VSS.n321 0.903568
R9193 VSS.n1223 VSS.n1219 0.903568
R9194 VSS.n1303 VSS.n1275 0.903568
R9195 VSS.n4051 VSS.n4010 0.903568
R9196 VSS.n3920 VSS.n3867 0.903568
R9197 VSS.n5412 VSS.n5411 0.871989
R9198 VSS.n130 VSS.n124 0.871989
R9199 VSS.n5405 VSS.n132 0.871989
R9200 VSS.n5404 VSS.n133 0.871989
R9201 VSS.n5389 VSS.n5388 0.871989
R9202 VSS.n5394 VSS.n5392 0.871989
R9203 VSS.n5393 VSS.n102 0.871989
R9204 VSS.n5418 VSS.n5417 0.871989
R9205 VSS.n5199 VSS.n5198 0.871989
R9206 VSS.n5168 VSS.n5160 0.871989
R9207 VSS.n5192 VSS.n5170 0.871989
R9208 VSS.n5191 VSS.n5171 0.871989
R9209 VSS.n5176 VSS.n5175 0.871989
R9210 VSS.n5181 VSS.n5179 0.871989
R9211 VSS.n5180 VSS.n401 0.871989
R9212 VSS.n5205 VSS.n5204 0.871989
R9213 VSS.n4946 VSS.n4945 0.871989
R9214 VSS.n4915 VSS.n4907 0.871989
R9215 VSS.n4939 VSS.n4917 0.871989
R9216 VSS.n4938 VSS.n4918 0.871989
R9217 VSS.n4923 VSS.n4922 0.871989
R9218 VSS.n4928 VSS.n4926 0.871989
R9219 VSS.n4927 VSS.n816 0.871989
R9220 VSS.n4952 VSS.n4951 0.871989
R9221 VSS.n3668 VSS.n3667 0.871989
R9222 VSS.n3632 VSS.n3624 0.871989
R9223 VSS.n3661 VSS.n3634 0.871989
R9224 VSS.n3660 VSS.n3635 0.871989
R9225 VSS.n3640 VSS.n3639 0.871989
R9226 VSS.n3650 VSS.n3643 0.871989
R9227 VSS.n3649 VSS.n3644 0.871989
R9228 VSS.n3646 VSS.n3645 0.871989
R9229 VSS.n5489 VSS.n53 0.871989
R9230 VSS.n5488 VSS.n54 0.871989
R9231 VSS.n5485 VSS.n50 0.871989
R9232 VSS.n49 VSS.n47 0.871989
R9233 VSS.n45 VSS.n44 0.871989
R9234 VSS.n5506 VSS.n40 0.871989
R9235 VSS.n5505 VSS.n41 0.871989
R9236 VSS.n5512 VSS.n36 0.871989
R9237 VSS.n4502 VSS.n70 0.82504
R9238 VSS.n966 VSS.n847 0.82504
R9239 VSS.n3680 VSS.n3478 0.82504
R9240 VSS.n5431 VSS.n83 0.82504
R9241 VSS.n4402 VSS.n1651 0.746512
R9242 VSS.n4991 VSS.n761 0.746512
R9243 VSS.n5231 VSS.n332 0.746512
R9244 VSS.n679 VSS.n321 0.746512
R9245 VSS.n1376 VSS.n1375 0.708416
R9246 VSS.n5401 VSS 0.599649
R9247 VSS.n5188 VSS 0.599649
R9248 VSS.n4935 VSS 0.599649
R9249 VSS.n3657 VSS 0.599649
R9250 VSS.n5498 VSS 0.599649
R9251 VSS.n1876 VSS.n1875 0.5301
R9252 VSS.n1877 VSS.n1876 0.5301
R9253 VSS.n4636 VSS.n4635 0.512067
R9254 VSS.n5348 VSS.n170 0.436245
R9255 VSS.n5345 VSS.n5344 0.436245
R9256 VSS.n182 VSS.n178 0.436245
R9257 VSS.n5338 VSS.n180 0.436245
R9258 VSS.n580 VSS.n573 0.436245
R9259 VSS.n584 VSS.n571 0.436245
R9260 VSS.n589 VSS.n587 0.436245
R9261 VSS.n594 VSS.n568 0.436245
R9262 VSS.n5328 VSS.n203 0.436245
R9263 VSS.n5325 VSS.n5324 0.436245
R9264 VSS.n223 VSS.n210 0.436245
R9265 VSS.n5318 VSS.n216 0.436245
R9266 VSS.n5313 VSS.n218 0.436245
R9267 VSS.n623 VSS.n622 0.436245
R9268 VSS.n632 VSS.n628 0.436245
R9269 VSS.n637 VSS.n614 0.436245
R9270 VSS.n5138 VSS.n424 0.436245
R9271 VSS.n5135 VSS.n5134 0.436245
R9272 VSS.n5130 VSS.n436 0.436245
R9273 VSS.n438 VSS.n437 0.436245
R9274 VSS.n858 VSS.n851 0.436245
R9275 VSS.n868 VSS.n865 0.436245
R9276 VSS.n872 VSS.n849 0.436245
R9277 VSS.n962 VSS.n874 0.436245
R9278 VSS.n4379 VSS.n1690 0.436245
R9279 VSS.n4376 VSS.n4375 0.436245
R9280 VSS.n1703 VSS.n1699 0.436245
R9281 VSS.n4369 VSS.n1701 0.436245
R9282 VSS.n1718 VSS.n1713 0.436245
R9283 VSS.n1728 VSS.n1725 0.436245
R9284 VSS.n1735 VSS.n1711 0.436245
R9285 VSS.n1737 VSS.n1407 0.436245
R9286 VSS.n4577 VSS.n4576 0.436245
R9287 VSS.n4572 VSS.n1448 0.436245
R9288 VSS.n4529 VSS.n1449 0.436245
R9289 VSS.n4566 VSS.n4563 0.436245
R9290 VSS.n4557 VSS.n4538 0.436245
R9291 VSS.n4543 VSS.n4539 0.436245
R9292 VSS.n4551 VSS.n4548 0.436245
R9293 VSS.n5532 VSS.n27 0.436245
R9294 VSS.n3674 VSS.n3481 0.436245
R9295 VSS.n3523 VSS.n3484 0.436245
R9296 VSS.n3528 VSS.n3527 0.436245
R9297 VSS.n3532 VSS.n3531 0.436245
R9298 VSS.n3559 VSS.n3517 0.436245
R9299 VSS.n3549 VSS.n3538 0.436245
R9300 VSS.n3546 VSS.n3545 0.436245
R9301 VSS.n1456 VSS.n1453 0.436245
R9302 VSS.n4493 VSS.n1476 0.436245
R9303 VSS.n4490 VSS.n4489 0.436245
R9304 VSS.n4485 VSS.n1487 0.436245
R9305 VSS.n1489 VSS.n1488 0.436245
R9306 VSS.n1635 VSS.n1626 0.436245
R9307 VSS.n1639 VSS.n1624 0.436245
R9308 VSS.n1644 VSS.n1622 0.436245
R9309 VSS.n1649 VSS.n1620 0.436245
R9310 VSS.n4885 VSS.n839 0.436245
R9311 VSS.n4882 VSS.n4881 0.436245
R9312 VSS.n4877 VSS.n974 0.436245
R9313 VSS.n976 VSS.n975 0.436245
R9314 VSS.n3464 VSS.n3463 0.436245
R9315 VSS.n3469 VSS.n3468 0.436245
R9316 VSS.n3473 VSS.n3472 0.436245
R9317 VSS.n3685 VSS.n3684 0.436245
R9318 VSS.n4866 VSS.n997 0.436245
R9319 VSS.n4863 VSS.n4862 0.436245
R9320 VSS.n4858 VSS.n1008 0.436245
R9321 VSS.n1010 VSS.n1009 0.436245
R9322 VSS.n3721 VSS.n3712 0.436245
R9323 VSS.n3725 VSS.n3710 0.436245
R9324 VSS.n3730 VSS.n3708 0.436245
R9325 VSS.n3735 VSS.n3706 0.436245
R9326 VSS.n5119 VSS.n459 0.436245
R9327 VSS.n5116 VSS.n5115 0.436245
R9328 VSS.n5111 VSS.n467 0.436245
R9329 VSS.n469 VSS.n468 0.436245
R9330 VSS.n926 VSS.n917 0.436245
R9331 VSS.n930 VSS.n915 0.436245
R9332 VSS.n935 VSS.n913 0.436245
R9333 VSS.n940 VSS.n911 0.436245
R9334 VSS.n3023 VSS.n3022 0.434398
R9335 VSS.n2858 VSS.n2857 0.434398
R9336 VSS.n3012 VSS.n2862 0.434398
R9337 VSS.n3008 VSS.n3007 0.434398
R9338 VSS.n2869 VSS.n2868 0.434398
R9339 VSS.n2998 VSS.n2873 0.434398
R9340 VSS.n2991 VSS.n2990 0.434398
R9341 VSS.n2986 VSS.n2878 0.434398
R9342 VSS.n2717 VSS.n2716 0.434398
R9343 VSS.n2081 VSS.n2080 0.434398
R9344 VSS.n2234 VSS.n2085 0.434398
R9345 VSS.n2230 VSS.n2229 0.434398
R9346 VSS.n2092 VSS.n2091 0.434398
R9347 VSS.n2220 VSS.n2096 0.434398
R9348 VSS.n2213 VSS.n2212 0.434398
R9349 VSS.n2208 VSS.n2207 0.434398
R9350 VSS.n3931 VSS.n3930 0.434398
R9351 VSS.n3281 VSS.n3280 0.434398
R9352 VSS.n3409 VSS.n3285 0.434398
R9353 VSS.n3405 VSS.n3404 0.434398
R9354 VSS.n3292 VSS.n3291 0.434398
R9355 VSS.n3395 VSS.n3296 0.434398
R9356 VSS.n3388 VSS.n3387 0.434398
R9357 VSS.n3383 VSS.n3301 0.434398
R9358 VSS.n4787 VSS.n1062 0.434398
R9359 VSS.n1064 VSS.n1063 0.434398
R9360 VSS.n4782 VSS.n1065 0.434398
R9361 VSS.n3843 VSS.n3835 0.434398
R9362 VSS.n3852 VSS.n3834 0.434398
R9363 VSS.n3856 VSS.n3833 0.434398
R9364 VSS.n3861 VSS.n3859 0.434398
R9365 VSS.n3865 VSS.n3831 0.434398
R9366 VSS.n4291 VSS.n1783 0.434398
R9367 VSS.n1785 VSS.n1784 0.434398
R9368 VSS.n4286 VSS.n1789 0.434398
R9369 VSS.n2465 VSS.n2458 0.434398
R9370 VSS.n2474 VSS.n2457 0.434398
R9371 VSS.n2478 VSS.n2454 0.434398
R9372 VSS.n2485 VSS.n2484 0.434398
R9373 VSS.n2489 VSS.n2488 0.434398
R9374 VSS.n2747 VSS.n2746 0.433481
R9375 VSS.n2742 VSS.n2068 0.433481
R9376 VSS.n2134 VSS.n2070 0.433481
R9377 VSS.n2136 VSS.n2127 0.433481
R9378 VSS.n2151 VSS.n2146 0.433481
R9379 VSS.n2149 VSS.n2124 0.433481
R9380 VSS.n2164 VSS.n2125 0.433481
R9381 VSS.n2161 VSS.n2160 0.433481
R9382 VSS.n3053 VSS.n3052 0.433481
R9383 VSS.n3048 VSS.n2025 0.433481
R9384 VSS.n2913 VSS.n2027 0.433481
R9385 VSS.n2915 VSS.n2906 0.433481
R9386 VSS.n2930 VSS.n2925 0.433481
R9387 VSS.n2928 VSS.n2903 0.433481
R9388 VSS.n2943 VSS.n2904 0.433481
R9389 VSS.n2940 VSS.n2939 0.433481
R9390 VSS.n4777 VSS.n1089 0.433481
R9391 VSS.n4759 VSS.n1093 0.433481
R9392 VSS.n1135 VSS.n1134 0.433481
R9393 VSS.n4754 VSS.n1136 0.433481
R9394 VSS.n4746 VSS.n1146 0.433481
R9395 VSS.n1150 VSS.n1149 0.433481
R9396 VSS.n4741 VSS.n1151 0.433481
R9397 VSS.n4738 VSS.n4737 0.433481
R9398 VSS.n3961 VSS.n3960 0.433481
R9399 VSS.n3956 VSS.n1949 0.433481
R9400 VSS.n3316 VSS.n1951 0.433481
R9401 VSS.n3318 VSS.n3309 0.433481
R9402 VSS.n3333 VSS.n3328 0.433481
R9403 VSS.n3331 VSS.n3307 0.433481
R9404 VSS.n3340 VSS.n3339 0.433481
R9405 VSS.n3967 VSS.n3966 0.433481
R9406 VSS.n1834 VSS.n1810 0.433481
R9407 VSS.n4278 VSS.n1811 0.433481
R9408 VSS.n1840 VSS.n1839 0.433481
R9409 VSS.n4246 VSS.n1842 0.433481
R9410 VSS.n4234 VSS.n1844 0.433481
R9411 VSS.n4229 VSS.n4226 0.433481
R9412 VSS.n4222 VSS.n1848 0.433481
R9413 VSS.n4220 VSS.n4217 0.433481
R9414 VSS.n5308 VSS.n242 0.433481
R9415 VSS.n5280 VSS.n246 0.433481
R9416 VSS.n273 VSS.n272 0.433481
R9417 VSS.n5275 VSS.n274 0.433481
R9418 VSS.n5267 VSS.n284 0.433481
R9419 VSS.n288 VSS.n287 0.433481
R9420 VSS.n5262 VSS.n289 0.433481
R9421 VSS.n5259 VSS.n5258 0.433481
R9422 VSS.n5101 VSS.n491 0.433481
R9423 VSS.n5073 VSS.n495 0.433481
R9424 VSS.n701 VSS.n700 0.433481
R9425 VSS.n5068 VSS.n702 0.433481
R9426 VSS.n5060 VSS.n712 0.433481
R9427 VSS.n716 VSS.n715 0.433481
R9428 VSS.n5055 VSS.n717 0.433481
R9429 VSS.n5052 VSS.n5051 0.433481
R9430 VSS.n4848 VSS.n1032 0.433481
R9431 VSS.n3777 VSS.n1036 0.433481
R9432 VSS.n3778 VSS.n3759 0.433481
R9433 VSS.n3783 VSS.n3758 0.433481
R9434 VSS.n3791 VSS.n3757 0.433481
R9435 VSS.n3794 VSS.n3756 0.433481
R9436 VSS.n3805 VSS.n3801 0.433481
R9437 VSS.n3810 VSS.n3754 0.433481
R9438 VSS.n4475 VSS.n1511 0.433481
R9439 VSS.n4447 VSS.n1515 0.433481
R9440 VSS.n1538 VSS.n1537 0.433481
R9441 VSS.n4442 VSS.n1539 0.433481
R9442 VSS.n4434 VSS.n1549 0.433481
R9443 VSS.n1553 VSS.n1552 0.433481
R9444 VSS.n4429 VSS.n1554 0.433481
R9445 VSS.n4426 VSS.n4425 0.433481
R9446 VSS.n4358 VSS.n1752 0.433481
R9447 VSS.n4355 VSS.n4354 0.433481
R9448 VSS.n4338 VSS.n1759 0.433481
R9449 VSS.n4348 VSS.n1761 0.433481
R9450 VSS.n2422 VSS.n2413 0.433481
R9451 VSS.n2427 VSS.n2412 0.433481
R9452 VSS.n2430 VSS.n2411 0.433481
R9453 VSS.n2511 VSS.n2510 0.433481
R9454 VSS.n1892 VSS.n1871 0.344944
R9455 VSS.n5333 VSS 0.300074
R9456 VSS VSS.n217 0.300074
R9457 VSS.n5125 VSS 0.300074
R9458 VSS.n4364 VSS 0.300074
R9459 VSS.n4535 VSS 0.300074
R9460 VSS.n3556 VSS 0.300074
R9461 VSS.n4480 VSS 0.300074
R9462 VSS.n4872 VSS 0.300074
R9463 VSS.n4853 VSS 0.300074
R9464 VSS.n5106 VSS 0.300074
R9465 VSS.n2993 VSS 0.298805
R9466 VSS.n2215 VSS 0.298805
R9467 VSS.n3390 VSS 0.298805
R9468 VSS.n3838 VSS 0.298805
R9469 VSS.n2460 VSS 0.298805
R9470 VSS.n2139 VSS 0.298174
R9471 VSS.n2918 VSS 0.298174
R9472 VSS.n4751 VSS 0.298174
R9473 VSS.n3321 VSS 0.298174
R9474 VSS.n4241 VSS 0.298174
R9475 VSS.n5272 VSS 0.298174
R9476 VSS.n5065 VSS 0.298174
R9477 VSS.n3786 VSS 0.298174
R9478 VSS.n4439 VSS 0.298174
R9479 VSS.n4343 VSS 0.298174
R9480 VSS VSS.n5400 0.27284
R9481 VSS VSS.n5187 0.27284
R9482 VSS VSS.n4934 0.27284
R9483 VSS VSS.n3656 0.27284
R9484 VSS VSS.n5497 0.27284
R9485 VSS.n1887 VSS.n1886 0.215691
R9486 VSS.n1894 VSS 0.140071
R9487 VSS.n575 VSS 0.13667
R9488 VSS.n616 VSS 0.13667
R9489 VSS.n857 VSS 0.13667
R9490 VSS.n1717 VSS 0.13667
R9491 VSS VSS.n4533 0.13667
R9492 VSS VSS.n3555 0.13667
R9493 VSS.n1630 VSS 0.13667
R9494 VSS.n3459 VSS 0.13667
R9495 VSS.n3716 VSS 0.13667
R9496 VSS.n921 VSS 0.13667
R9497 VSS.n3003 VSS 0.136093
R9498 VSS.n2225 VSS 0.136093
R9499 VSS.n3400 VSS 0.136093
R9500 VSS.n3847 VSS 0.136093
R9501 VSS.n2469 VSS 0.136093
R9502 VSS.n2128 VSS 0.135807
R9503 VSS.n2907 VSS 0.135807
R9504 VSS VSS.n4750 0.135807
R9505 VSS.n3310 VSS 0.135807
R9506 VSS VSS.n4238 0.135807
R9507 VSS VSS.n5271 0.135807
R9508 VSS VSS.n5064 0.135807
R9509 VSS.n3765 VSS 0.135807
R9510 VSS VSS.n4438 0.135807
R9511 VSS.n2421 VSS 0.135807
R9512 VSS.n1892 VSS 0.0664299
R9513 VSS.n5400 VSS 0.0549681
R9514 VSS.n5187 VSS 0.0549681
R9515 VSS.n4934 VSS 0.0549681
R9516 VSS.n3656 VSS 0.0549681
R9517 VSS.n5497 VSS 0.0549681
R9518 VSS.n4630 VSS.n1398 0.0338012
R9519 VSS.n1894 VSS.n1893 0.0280822
R9520 VSS.n2299 VSS.n2277 0.027734
R9521 VSS VSS.n575 0.027734
R9522 VSS.n2357 VSS.n2356 0.027734
R9523 VSS.n616 VSS 0.027734
R9524 VSS VSS.n857 0.027734
R9525 VSS VSS.n1717 0.027734
R9526 VSS VSS.n4533 0.027734
R9527 VSS.n3555 VSS 0.027734
R9528 VSS VSS.n1630 0.027734
R9529 VSS VSS.n3459 0.027734
R9530 VSS VSS.n3716 0.027734
R9531 VSS VSS.n921 0.027734
R9532 VSS.n3003 VSS 0.0276186
R9533 VSS.n2225 VSS 0.0276186
R9534 VSS.n3400 VSS 0.0276186
R9535 VSS VSS.n3847 0.0276186
R9536 VSS VSS.n2469 0.0276186
R9537 VSS.n4631 VSS.n1396 0.0275781
R9538 VSS.n2684 VSS.n2683 0.0275613
R9539 VSS.n2128 VSS 0.0275613
R9540 VSS.n2907 VSS 0.0275613
R9541 VSS.n4750 VSS 0.0275613
R9542 VSS.n3310 VSS 0.0275613
R9543 VSS.n4238 VSS 0.0275613
R9544 VSS.n4212 VSS.n4211 0.0275613
R9545 VSS.n2251 VSS.n267 0.0275613
R9546 VSS.n5271 VSS 0.0275613
R9547 VSS.n5064 VSS 0.0275613
R9548 VSS.n3765 VSS 0.0275613
R9549 VSS.n4438 VSS 0.0275613
R9550 VSS VSS.n2421 0.0275613
R9551 VSS.n2531 VSS.n2516 0.0275613
R9552 VSS VSS.n1882 0.0207703
R9553 VSS.n1879 VSS.n1878 0.0183341
R9554 VSS.n1888 VSS.n1887 0.0114834
R9555 VSS.n1878 VSS 0.00825612
R9556 VSS.n1895 VSS.n1892 0.00600823
R9557 VSS.n4636 VSS.n0 0.00569031
R9558 VSS.n1880 VSS.n1879 0.00459091
R9559 VSS.n1895 VSS.n1894 0.00399193
R9560 VSS.n4633 VSS.n4632 0.00134175
R9561 VSS.n1888 VSS 0.00123972
R9562 MINUS.n6 MINUS.n5 280.983
R9563 MINUS.n1 MINUS.n0 83.5719
R9564 MINUS.n11 MINUS.n10 83.5719
R9565 MINUS.n14 MINUS.n1 73.8498
R9566 MINUS.n4 MINUS.t4 67.4224
R9567 MINUS.n4 MINUS.t5 66.2083
R9568 MINUS.t3 MINUS.n9 64.5544
R9569 MINUS.n10 MINUS.n1 26.074
R9570 MINUS.n7 MINUS.t0 11.6945
R9571 MINUS MINUS.n4 11.4492
R9572 MINUS.n8 MINUS.n7 3.79884
R9573 MINUS.n5 MINUS.t1 2.857
R9574 MINUS.n5 MINUS.t2 2.857
R9575 MINUS.n6 MINUS 2.00148
R9576 MINUS.n13 MINUS.n12 1.5505
R9577 MINUS.n3 MINUS.n2 1.5505
R9578 MINUS.n9 MINUS.n8 1.49631
R9579 MINUS.n9 MINUS.n3 1.41981
R9580 MINUS.n11 MINUS.n3 1.07024
R9581 MINUS.n12 MINUS.n0 0.885803
R9582 MINUS.n12 MINUS.n11 0.77514
R9583 MINUS MINUS.n0 0.756696
R9584 MINUS.n14 MINUS.n13 0.71401
R9585 MINUS MINUS.n14 0.576402
R9586 MINUS.n10 MINUS.t3 0.290206
R9587 MINUS.n13 MINUS.n2 0.0205321
R9588 MINUS.n7 MINUS.n6 0.00659756
R9589 MINUS.n8 MINUS.n2 0.00130128
R9590 a_17692_n8717.n0 a_17692_n8717.n3 215.76
R9591 a_17692_n8717.n0 a_17692_n8717.n2 215
R9592 a_17692_n8717.n1 a_17692_n8717.t9 192.987
R9593 a_17692_n8717.n1 a_17692_n8717.t8 192.987
R9594 a_17692_n8717.n1 a_17692_n8717.t2 192.475
R9595 a_17692_n8717.n1 a_17692_n8717.t4 192.475
R9596 a_17692_n8717.n4 a_17692_n8717.n0 154.554
R9597 a_17692_n8717.t5 a_17692_n8717.n4 7.14175
R9598 a_17692_n8717.n4 a_17692_n8717.t3 7.14175
R9599 a_17692_n8717.n0 a_17692_n8717.n1 6.97315
R9600 a_17692_n8717.n3 a_17692_n8717.t6 2.1755
R9601 a_17692_n8717.n3 a_17692_n8717.t0 2.1755
R9602 a_17692_n8717.n2 a_17692_n8717.t1 2.1755
R9603 a_17692_n8717.n2 a_17692_n8717.t7 2.1755
R9604 Vbgr.n1 Vbgr.n0 275.454
R9605 Vbgr Vbgr.t0 23.4071
R9606 Vbgr.n5 Vbgr.n1 8.18097
R9607 Vbgr.n2 Vbgr.t5 4.9747
R9608 Vbgr.n4 Vbgr.t4 4.91993
R9609 Vbgr.n3 Vbgr.t3 4.91993
R9610 Vbgr.n2 Vbgr.t6 4.91993
R9611 Vbgr.n1 Vbgr 3.01173
R9612 Vbgr.n0 Vbgr.t2 2.857
R9613 Vbgr.n0 Vbgr.t1 2.857
R9614 Vbgr Vbgr.n4 2.30408
R9615 Vbgr Vbgr.n5 0.0633049
R9616 Vbgr.n5 Vbgr 0.0626981
R9617 Vbgr.n4 Vbgr.n3 0.0552707
R9618 Vbgr.n3 Vbgr.n2 0.0552707
R9619 Sop.n2 Sop.n1 210.935
R9620 Sop.n2 Sop.n0 210.935
R9621 Sop Sop.n3 78.6661
R9622 Sop.n3 Sop.t0 8.7005
R9623 Sop.n3 Sop.t1 8.7005
R9624 Sop Sop.n2 5.60828
R9625 Sop.n0 Sop.t5 2.1755
R9626 Sop.n0 Sop.t3 2.1755
R9627 Sop.n1 Sop.t2 2.1755
R9628 Sop.n1 Sop.t4 2.1755
C0 a_24244_n9724# a_24323_n8877# 0.033727f
C1 Vbgr a_25579_n8877# 0.030096f
C2 a_25081_n8277# a_23991_n8277# 0.340116f
C3 a_24478_n10376# a_25414_n10376# 4.82e-21
C4 a_24946_n10376# a_25180_n9724# 0.034607f
C5 a_23493_n8277# a_23659_n8877# 0.023433f
C6 MINUS a_25180_n9724# 0.009501f
C7 MINUS a_25247_n8277# 0.152215f
C8 Vbgr a_24323_n8877# 2.61e-19
C9 XQ2[0|0].Emitter a_24712_n9724# 0.059011f
C10 XQ2[0|0].Emitter a_24915_n8877# 0.112162f
C11 MINUS a_23659_n8877# 0.001756f
C12 Vbgr a_24244_n9724# 1.56e-20
C13 a_23659_n8877# a_23991_n8277# 0.003644f
C14 a_24010_n10376# a_24478_n10376# 0.298666f
C15 VDD MINUS 1.06539f
C16 a_24712_n9724# a_24323_n8877# 0.042461f
C17 XQ2[0|0].Emitter a_24946_n10376# 0.003391f
C18 MINUS a_23825_n8877# 0.001691f
C19 a_24915_n8877# a_24323_n8877# 0.453352f
C20 a_24010_n10376# a_23776_n9724# 0.034605f
C21 MINUS XQ2[0|0].Emitter 4.67044f
C22 a_25180_n9724# a_25414_n10376# 0.034603f
C23 VDD a_23991_n8277# 4.51e-19
C24 MINUS a_25579_n8877# 0.394455f
C25 a_23659_n8877# a_24157_n8277# 0.023451f
C26 a_23825_n8877# a_23991_n8277# 0.023433f
C27 a_24244_n9724# a_24712_n9724# 0.298808f
C28 XQ2[0|0].Emitter a_23991_n8277# 0.001537f
C29 a_24946_n10376# a_24323_n8877# 0.004947f
C30 Gcm2 Sop 0.116649f
C31 MINUS a_24323_n8877# 0.355534f
C32 Vbgr a_24712_n9724# 1.13e-19
C33 VDD a_24157_n8277# 9.21e-19
C34 a_23991_n8277# a_24323_n8877# 0.017118f
C35 XQ2[0|0].Emitter a_25414_n10376# 0.003384f
C36 Vbgr a_23493_n8277# 1.82e-19
C37 a_25579_n8877# a_25414_n10376# 0.002985f
C38 a_24010_n10376# a_23659_n8877# 0.003748f
C39 Vbgr MINUS 0.420749f
C40 a_24157_n8277# a_24323_n8877# 0.023433f
C41 a_23542_n10376# a_24946_n10376# 3.11e-21
C42 a_24244_n9724# a_24157_n8277# 0.002284f
C43 a_24712_n9724# a_24946_n10376# 0.034601f
C44 MINUS a_24915_n8877# 0.006395f
C45 Vbgr a_25414_n10376# 0.033913f
C46 VDD Sop 0.021357f
C47 MINUS a_23493_n8277# 0.007454f
C48 a_24915_n8877# a_23991_n8277# 0.023915f
C49 a_23659_n8877# a_23776_n9724# 0.042257f
C50 a_25081_n8277# a_25180_n9724# 0.001698f
C51 a_25081_n8277# a_25247_n8277# 0.737085f
C52 VDD Gcm2 1.06632f
C53 a_23493_n8277# a_23991_n8277# 1.41e-19
C54 a_23542_n10376# a_25414_n10376# 6.09e-22
C55 a_24010_n10376# a_24244_n9724# 0.034611f
C56 Gcm2 a_23825_n8877# 0.002409f
C57 XQ2[0|0].Emitter a_24478_n10376# 0.002121f
C58 Gcm2 XQ2[0|0].Emitter 1.34e-19
C59 MINUS a_23991_n8277# 0.026436f
C60 a_25247_n8277# a_25180_n9724# 0.003106f
C61 VDD a_25081_n8277# 1.37e-19
C62 a_24478_n10376# a_24323_n8877# 0.004861f
C63 XQ2[0|0].Emitter a_25081_n8277# 0.001639f
C64 a_24010_n10376# a_23542_n10376# 0.298736f
C65 MINUS a_24157_n8277# 0.004856f
C66 a_24946_n10376# a_25414_n10376# 0.299281f
C67 a_25081_n8277# a_25579_n8877# 0.023915f
C68 a_24244_n9724# a_24478_n10376# 0.034612f
C69 a_23991_n8277# a_24157_n8277# 0.432514f
C70 XQ2[0|0].Emitter a_25180_n9724# 0.058405f
C71 XQ2[0|0].Emitter a_25247_n8277# 9.32e-19
C72 a_24244_n9724# a_23776_n9724# 0.298213f
C73 a_25081_n8277# a_24323_n8877# 0.003676f
C74 Vbgr Gcm2 0.006361f
C75 a_23659_n8877# a_23825_n8877# 0.745688f
C76 XQ2[0|0].Emitter a_23659_n8877# 0.004761f
C77 Vbgr a_23776_n9724# 3.15e-21
C78 a_25180_n9724# a_24323_n8877# 0.015496f
C79 a_25247_n8277# a_24323_n8877# 0.023915f
C80 a_24478_n10376# a_23542_n10376# 7.87e-20
C81 VDD XQ2[0|0].Emitter 0.264496f
C82 XQ2[0|0].Emitter a_23825_n8877# 0.002687f
C83 a_23542_n10376# a_23776_n9724# 0.034723f
C84 a_23659_n8877# a_24323_n8877# 0.337637f
C85 a_24478_n10376# a_24712_n9724# 0.034601f
C86 XQ2[0|0].Emitter a_25579_n8877# 0.024517f
C87 MINUS Sop 3.07732f
C88 Gcm2 a_23493_n8277# 0.016232f
C89 Vbgr a_25180_n9724# 0.297712f
C90 XQ2[0|0].Emitter a_24323_n8877# 0.381626f
C91 a_24478_n10376# a_24946_n10376# 0.298765f
C92 a_24010_n10376# a_25414_n10376# 1.89e-21
C93 Gcm2 MINUS 0.394647f
C94 a_24915_n8877# a_25081_n8277# 0.023915f
C95 a_25579_n8877# a_24323_n8877# 0.001551f
C96 Gcm2 a_23991_n8277# 0.078689f
C97 a_24712_n9724# a_25180_n9724# 0.29801f
C98 a_23659_n8877# a_23542_n10376# 0.004809f
C99 VDD Vbgr 3.54031f
C100 MINUS a_25081_n8277# 0.151236f
C101 Vbgr XQ2[0|0].Emitter 0.744237f
C102 Vbgr VSS 13.140335f
C103 VDD VSS 35.164814f
C104 a_25414_n10376# VSS 0.806369f
C105 a_25180_n9724# VSS 0.467234f
C106 a_24946_n10376# VSS 0.505692f
C107 a_24712_n9724# VSS 0.462354f
C108 a_24478_n10376# VSS 0.505614f
C109 a_24244_n9724# VSS 0.466284f
C110 a_24010_n10376# VSS 0.506957f
C111 a_23776_n9724# VSS 0.754256f
C112 a_23542_n10376# VSS 0.837674f
C113 a_25579_n8877# VSS 0.639712f
C114 a_25247_n8277# VSS 0.315247f
C115 a_25081_n8277# VSS 0.444742f
C116 a_24915_n8877# VSS 0.476392f
C117 a_24323_n8877# VSS 0.820643f
C118 a_24157_n8277# VSS 0.450227f
C119 a_23991_n8277# VSS 1.18248f
C120 a_23825_n8877# VSS 0.336082f
C121 a_23659_n8877# VSS 0.815395f
C122 a_23493_n8277# VSS 0.987762f
C123 Sop VSS 1.848726f
C124 XQ2[0|0].Emitter VSS 77.892204f
C125 MINUS VSS 7.369028f
C126 Gcm2 VSS 5.03475f
C127 Sop.t5 VSS 0.027992f
C128 Sop.t3 VSS 0.027992f
C129 Sop.n0 VSS 0.09895f
C130 Sop.t2 VSS 0.027992f
C131 Sop.t4 VSS 0.027992f
C132 Sop.n1 VSS 0.098958f
C133 Sop.n2 VSS 2.64181f
C134 Sop.t0 VSS 0.006998f
C135 Sop.t1 VSS 0.006998f
C136 Sop.n3 VSS 0.020916f
C137 Vbgr.t0 VSS 0.065722f
C138 Vbgr.t2 VSS 0.047673f
C139 Vbgr.t1 VSS 0.047673f
C140 Vbgr.n0 VSS 0.164993f
C141 Vbgr.n1 VSS 0.88215f
C142 Vbgr.t5 VSS 1.02041f
C143 Vbgr.t6 VSS 1.00728f
C144 Vbgr.n2 VSS 2.41934f
C145 Vbgr.t3 VSS 1.00728f
C146 Vbgr.n3 VSS 1.23703f
C147 Vbgr.t4 VSS 1.00728f
C148 Vbgr.n4 VSS 1.23062f
C149 Vbgr.n5 VSS 0.853808f
C150 a_17692_n8717.n0 VSS 1.2128f
C151 a_17692_n8717.n1 VSS 0.347951f
C152 a_17692_n8717.t3 VSS 0.018559f
C153 a_17692_n8717.t8 VSS 0.229926f
C154 a_17692_n8717.t4 VSS 0.229705f
C155 a_17692_n8717.t9 VSS 0.229926f
C156 a_17692_n8717.t2 VSS 0.229705f
C157 a_17692_n8717.t1 VSS 0.037118f
C158 a_17692_n8717.t7 VSS 0.037118f
C159 a_17692_n8717.n2 VSS 0.13831f
C160 a_17692_n8717.t6 VSS 0.037118f
C161 a_17692_n8717.t0 VSS 0.037118f
C162 a_17692_n8717.n3 VSS 0.139247f
C163 a_17692_n8717.n4 VSS 0.056842f
C164 a_17692_n8717.t5 VSS 0.018559f
C165 MINUS.n0 VSS 0.054958f
C166 MINUS.n1 VSS 0.249114f
C167 MINUS.n2 VSS 0.057743f
C168 MINUS.n3 VSS 0.102688f
C169 MINUS.t5 VSS 1.85662f
C170 MINUS.t4 VSS 1.86887f
C171 MINUS.n4 VSS 1.55839f
C172 MINUS.t1 VSS 0.051607f
C173 MINUS.t2 VSS 0.051607f
C174 MINUS.n5 VSS 0.184016f
C175 MINUS.n6 VSS 0.435286f
C176 MINUS.t0 VSS 0.172289f
C177 MINUS.n7 VSS 0.860588f
C178 MINUS.n8 VSS 1.31424f
C179 MINUS.n9 VSS 0.291197f
C180 MINUS.t3 VSS 0.204f
C181 MINUS.n10 VSS 0.055059f
C182 MINUS.n11 VSS 0.061751f
C183 MINUS.n12 VSS 0.055575f
C184 MINUS.n13 VSS 0.412266f
C185 MINUS.n14 VSS 0.281274f
C186 VDD.t33 VSS 0.255619f
C187 VDD.t29 VSS 0.042188f
C188 VDD.n0 VSS 0.068489f
C189 VDD.t18 VSS 0.311083f
C190 VDD.t31 VSS 0.444189f
C191 VDD.t27 VSS 0.107724f
C192 VDD.n1 VSS 0.093858f
C193 VDD.t1 VSS 0.008704f
C194 VDD.t36 VSS 0.008704f
C195 VDD.n2 VSS 0.026355f
C196 VDD.n3 VSS 0.1042f
C197 VDD.t19 VSS 0.008704f
C198 VDD.t34 VSS 0.008704f
C199 VDD.n4 VSS 0.026355f
C200 VDD.n5 VSS 0.1042f
C201 VDD.t30 VSS 0.107724f
C202 VDD.n6 VSS 0.093858f
C203 VDD.t32 VSS 0.042188f
C204 VDD.n7 VSS 0.065415f
C205 VDD.n8 VSS 0.562605f
C206 VDD.n9 VSS 0.099834f
C207 VDD.n10 VSS 0.18956f
C208 VDD.t24 VSS 0.123264f
C209 VDD.n11 VSS 0.09873f
C210 VDD.t20 VSS 0.123225f
C211 VDD.t26 VSS 0.139592f
C212 VDD.t11 VSS 0.021759f
C213 VDD.n12 VSS 0.075291f
C214 VDD.n13 VSS 0.092282f
C215 VDD.t3 VSS 0.021759f
C216 VDD.t7 VSS 0.021759f
C217 VDD.n14 VSS 0.075291f
C218 VDD.n15 VSS 0.086431f
C219 VDD.t13 VSS 0.021759f
C220 VDD.t17 VSS 0.021759f
C221 VDD.n16 VSS 0.075291f
C222 VDD.n17 VSS 0.086431f
C223 VDD.t5 VSS 0.021759f
C224 VDD.t9 VSS 0.021759f
C225 VDD.n18 VSS 0.075291f
C226 VDD.n19 VSS 0.086431f
C227 VDD.t15 VSS 0.021759f
C228 VDD.t22 VSS 0.021759f
C229 VDD.n20 VSS 0.075291f
C230 VDD.n21 VSS 0.093295f
C231 VDD.n22 VSS 0.099754f
C232 VDD.n23 VSS 0.047614f
C233 VDD.t23 VSS 0.117834f
C234 VDD.n24 VSS 0.191364f
C235 VDD.n25 VSS 0.476249f
C236 VDD.t21 VSS 0.423597f
C237 VDD.t14 VSS 0.256303f
C238 VDD.t8 VSS 0.256303f
C239 VDD.t4 VSS 0.256303f
C240 VDD.t16 VSS 0.256303f
C241 VDD.t12 VSS 0.256303f
C242 VDD.t6 VSS 0.256303f
C243 VDD.t2 VSS 0.256303f
C244 VDD.t10 VSS 0.256303f
C245 VDD.t25 VSS 0.401471f
C246 VDD.n26 VSS 0.316901f
C247 VDD.n27 VSS 0.04885f
C248 VDD.n28 VSS 0.210599f
C249 VDD.n29 VSS 0.434057f
C250 VDD.n30 VSS 0.257869f
C251 VDD.n31 VSS 0.014124f
C252 VDD.n32 VSS 0.504599f
C253 VDD.n33 VSS 0.596912f
C254 VDD.t28 VSS 0.450855f
C255 VDD.t35 VSS 0.311083f
C256 VDD.t0 VSS 0.211006f
C257 a_17750_n8805.t2 VSS 0.021553f
C258 a_17750_n8805.t1 VSS 0.021553f
C259 a_17750_n8805.n0 VSS 0.074808f
C260 a_17750_n8805.t5 VSS 0.775365f
C261 a_17750_n8805.t4 VSS 0.789346f
C262 a_17750_n8805.n1 VSS 0.997031f
C263 a_17750_n8805.n2 VSS 0.344677f
C264 a_17750_n8805.t3 VSS 0.025867f
C265 a_17750_n8805.n3 VSS 0.239533f
C266 a_17750_n8805.t0 VSS 0.010265f
C267 w_21453_n6696.t4 VSS 0.190494f
C268 w_21453_n6696.n0 VSS 2.8056f
C269 w_21453_n6696.n1 VSS 0.93363f
C270 w_21453_n6696.t3 VSS 0.017238f
C271 w_21453_n6696.t8 VSS 0.017238f
C272 w_21453_n6696.t5 VSS 0.017238f
C273 w_21453_n6696.n2 VSS 0.052919f
C274 w_21453_n6696.t16 VSS 0.243964f
C275 w_21453_n6696.t20 VSS 0.243954f
C276 w_21453_n6696.t18 VSS 0.243954f
C277 w_21453_n6696.t15 VSS 0.243954f
C278 w_21453_n6696.t13 VSS 0.243954f
C279 w_21453_n6696.t19 VSS 0.243954f
C280 w_21453_n6696.t17 VSS 0.243954f
C281 w_21453_n6696.t14 VSS 0.243954f
C282 w_21453_n6696.t2 VSS 0.015834f
C283 w_21453_n6696.t7 VSS 0.015834f
C284 w_21453_n6696.t1 VSS 1.9088f
C285 w_21453_n6696.t6 VSS 1.16234f
C286 w_21453_n6696.t9 VSS 1.9088f
C287 w_21453_n6696.t11 VSS 1.16234f
C288 w_21453_n6696.n3 VSS 1.03881f
C289 w_21453_n6696.t12 VSS 0.015834f
C290 w_21453_n6696.t10 VSS 0.015834f
C291 w_21453_n6696.n4 VSS 0.052329f
C292 w_21453_n6696.t0 VSS 0.017238f
.ends

