** sch_path: /home/ttuser/tt08-bgr/xschem/core_PreL.sch
.subckt core_PreL MINUS PLUS Vbgr VDD VSS vp
*.PININFO MINUS:O PLUS:O Vbgr:O VDD:I VSS:I vp:I
XQ1 VSS VSS MINUS sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
XQ2 VSS VSS net1 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=29
XM1 MINUS vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XM2 PLUS vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XM3 Vbgr vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XR19 net1 PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=0.93 mult=1 m=1
XR2 VSS PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6.35 mult=1 m=1
XR3 VSS MINUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6.35 mult=1 m=1
XR1 VSS Vbgr VSS sky130_fd_pr__res_xhigh_po_1p41 L=26.57 mult=1 m=1
.ends
.end
