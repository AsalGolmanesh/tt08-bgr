** sch_path: /home/ttuser/tt08-bgr/xschem/BGRwOpampRes.sch
**.subckt BGRwOpampRes
XQ1 VSS VSS MINUS sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ2 VSS VSS net8 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=33
XM1 net1 vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vbgr vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 VDD GND 1.8
V2 VSS GND 0
Vmeas net1 MINUS 0
.save i(vmeas)
Vmeas1 net2 PLUS 0
.save i(vmeas1)
.save v(vdd)
.save v(net1)
.save v(vdd)
.save v(net2)
.save v(vdd)
.save v(vbgr)
XM4 vp MINUS net3 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net5 PLUS net3 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 vp net5 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.save v(vp)
.save v(net3)
.save v(net5)
.save v(net3)
XM10 net6 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net5 net5 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.save v(vdd)
.save v(net5)
.save v(vdd)
.save v(vp)
.save v(net6)
.save v(vss)
.save v(net4)
.save v(vss)
Vmeas3 net3 net6 0
.save i(vmeas3)
XM8 net7 vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas2 net7 net4 0
.save i(vmeas2)
.save v(vdd)
.save v(net7)
XR2 VSS PLUS VSS sky130_fd_pr__res_xhigh_po W=1 L=22 mult=1 m=1
XR3 VSS MINUS VSS sky130_fd_pr__res_xhigh_po W=1 L=22 mult=1 m=1
XM11 VSS Vbgr vp vp sky130_fd_pr__pfet_01v8_lvt L=1 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.save v(minus)
.save v(plus)
XR28 net8 PLUS VSS sky130_fd_pr__res_xhigh_po W=1 L=4 mult=1 m=1
XR1 VSS Vbgr VSS sky130_fd_pr__res_xhigh_po W=1 L=24 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
**** begin user architecture code



.options savecurrents
.control


save @m.xm1.msky130_fd_pr__ppet_01v8_lvt[gm]
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[vgs]
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[cgg]
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm1.msky130_fd_pr__pfet_01v8_lvt[vth]


save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vgs]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[cgg]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm2.msky130_fd_pr__pfet_01v8_lvt[vth]


save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[vgs]
save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[cgg]
save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[vth]

save @q.xq1.qsky130_fd_pr__pnp_05v5_W3p40L3p40[vbe]
save @q.xq2.qsky130_fd_pr__pnp_05v5_W3p40L3p40[vbe]


save @m.xm6.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm6.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vgs]
save @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm6.msky130_fd_pr__pfet_01v8_lvt[cgg]
save @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vth]

save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[vgs]
save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[cgg]
save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm7.msky130_fd_pr__pfet_01v8_lvt[vth]



save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[gm]
save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[id]
save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[vgs]
save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[vds]
save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[cgg]
save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[vdsat]
save @m.xm8.msky130_fd_pr__pfet_01v8_lvt[vth]


save @m.xm4.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm4.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vgs]
save @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm4.msky130_fd_pr__nfet_01v8_lvt[cgg]
save @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vth]


save @m.xm5.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm5.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm5.msky130_fd_pr__nfet_01v8_lvt[vgs]
save @m.xm5.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm5.msky130_fd_pr__nfet_01v8_lvt[cgg]
save @m.xm5.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm5.msky130_fd_pr__nfet_01v8_lvt[vth]



save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[vgs]
save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[cgg]
save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[vth]



save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[vgs]
save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[cgg]
save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[vth]


save @m.xm11.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm11.msky130_fd_pr__nfet_01v8_lvt[id]
save @m.xm11.msky130_fd_pr__nfet_01v8_lvt[vgs]
save @m.xm11.msky130_fd_pr__nfet_01v8_lvt[vds]
save @m.xm11.msky130_fd_pr__nfet_01v8_lvt[cgg]
save @m.xm11.msky130_fd_pr__nfet_01v8_lvt[vdsat]
save @m.xm11.msky130_fd_pr__nfet_01v8_lvt[vth]
save all
op
write BGRwOpampRes.raw
dc TEMP -40 125 10
plot Vbgr
*tran 20p 2u
*write BGRwOpampRes_startup.raw
.endc



**** end user architecture code
.end
