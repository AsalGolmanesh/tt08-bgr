magic
tech sky130A
magscale 1 2
timestamp 1725319194
<< nwell >>
rect 24100 -4757 24530 -4756
rect 18142 -6992 20748 -5385
rect 24100 -6921 24702 -4757
rect 26205 -6494 26499 -4753
rect 26188 -6918 26499 -6494
<< pwell >>
rect 23255 -7850 23397 -7798
rect 23991 -7845 24061 -7746
rect 25081 -7845 25151 -7739
rect 25745 -7873 25815 -7823
rect 25911 -7856 26147 -7832
rect 26054 -7995 26115 -7856
rect 23178 -8122 23243 -8091
rect 23247 -8878 23297 -8621
rect 26054 -8685 26138 -7995
rect 25413 -8868 25538 -8863
rect 24323 -8978 24393 -8877
rect 25413 -8953 25550 -8868
rect 26054 -8874 26115 -8685
rect 25911 -8910 26147 -8874
rect 25413 -8978 25483 -8953
rect 25490 -8955 25550 -8953
rect 26155 -9258 26179 -9227
rect 23165 -9708 23444 -9297
rect 25775 -9360 25776 -9260
rect 25891 -9394 26179 -9258
rect 23167 -9808 23234 -9708
rect 26155 -9947 26179 -9394
rect 23212 -10359 23433 -9964
rect 25889 -10512 26149 -10332
<< nbase >>
rect 29575 -9292 29614 -9291
<< pdiff >>
rect 29575 -9292 29614 -9291
<< psubdiff >>
rect 16171 -3802 16195 -3600
rect 33602 -3802 33626 -3600
rect 16200 -4004 16402 -3980
rect 33402 -4202 33606 -4178
rect 16539 -7193 16714 -7082
rect 16539 -8666 16594 -7193
rect 16686 -8666 16714 -7193
rect 16539 -8795 16714 -8666
rect 22099 -7202 22274 -7091
rect 22099 -8675 22154 -7202
rect 22246 -8675 22274 -7202
rect 22099 -8804 22274 -8675
rect 18765 -9426 18971 -9399
rect 18765 -9787 18825 -9426
rect 18890 -9787 18971 -9426
rect 18765 -9800 18971 -9787
rect 20067 -9421 20272 -9394
rect 20067 -9782 20126 -9421
rect 20191 -9782 20272 -9421
rect 20067 -9795 20272 -9782
rect 33402 -12426 33606 -12402
rect 16200 -12624 16402 -12600
rect 16172 -12997 16196 -12799
rect 33598 -12997 33622 -12799
<< nsubdiff >>
rect 24300 -4967 24403 -4901
rect 18263 -5747 18531 -5684
rect 18263 -6691 18321 -5747
rect 18455 -6691 18531 -5747
rect 18263 -6806 18531 -6691
rect 20334 -5734 20602 -5671
rect 20334 -6678 20392 -5734
rect 20526 -6678 20602 -5734
rect 20334 -6793 20602 -6678
rect 24300 -6747 24329 -4967
rect 24372 -6747 24403 -4967
rect 24300 -6802 24403 -6747
rect 26305 -4967 26408 -4901
rect 26305 -6747 26334 -4967
rect 26377 -6747 26408 -4967
rect 26305 -6802 26408 -6747
<< psubdiffcont >>
rect 16195 -3802 33602 -3600
rect 16200 -12600 16402 -4004
rect 16594 -8666 16686 -7193
rect 22154 -8675 22246 -7202
rect 18825 -9787 18890 -9426
rect 20126 -9782 20191 -9421
rect 33402 -12402 33606 -4202
rect 16196 -12997 33598 -12799
<< nsubdiffcont >>
rect 18321 -6691 18455 -5747
rect 20392 -6678 20526 -5734
rect 24329 -6747 24372 -4967
rect 26334 -6747 26377 -4967
<< locali >>
rect 16179 -3802 16195 -3600
rect 33602 -3802 33618 -3600
rect 16202 -3988 16402 -3802
rect 16200 -4004 16402 -3988
rect 33400 -4100 33602 -3802
rect 33400 -4174 33606 -4100
rect 33402 -4202 33606 -4174
rect 26630 -4488 33006 -4471
rect 26630 -4707 33070 -4488
rect 18289 -5747 18487 -5726
rect 18289 -6069 18320 -5747
rect 18289 -6691 18321 -6069
rect 18455 -6691 18487 -5747
rect 18289 -6745 18487 -6691
rect 20360 -5734 20558 -5713
rect 20360 -6678 20392 -5734
rect 20526 -5735 20558 -5734
rect 20528 -6067 20558 -5735
rect 20526 -6678 20558 -6067
rect 24317 -6221 24329 -5200
rect 24372 -6221 24384 -5200
rect 20360 -6732 20558 -6678
rect 24317 -6720 24319 -6221
rect 26322 -6225 26334 -5200
rect 26377 -6225 26389 -5200
rect 26631 -5996 33071 -5523
rect 24317 -6747 24329 -6720
rect 24372 -6747 24384 -6720
rect 24317 -6784 24384 -6747
rect 26322 -6747 26334 -6724
rect 26377 -6747 26389 -6724
rect 26322 -6784 26389 -6747
rect 16571 -7193 16700 -7119
rect 16402 -7774 16405 -7506
rect 16571 -8116 16594 -7193
rect 16686 -8116 16700 -7193
rect 16571 -8665 16591 -8116
rect 16687 -8665 16700 -8116
rect 16571 -8666 16594 -8665
rect 16686 -8666 16700 -8665
rect 16571 -8772 16700 -8666
rect 22131 -7202 22260 -7128
rect 22131 -8125 22154 -7202
rect 22246 -8125 22260 -7202
rect 26630 -7284 33073 -6813
rect 22131 -8674 22151 -8125
rect 22247 -8674 22260 -8125
rect 26627 -8572 33072 -8099
rect 22131 -8675 22154 -8674
rect 22246 -8675 22260 -8674
rect 22131 -8781 22260 -8675
rect 29575 -9292 29614 -9291
rect 18809 -9426 18915 -9401
rect 18809 -9787 18825 -9426
rect 18890 -9787 18915 -9426
rect 18809 -9804 18915 -9787
rect 20110 -9421 20216 -9396
rect 20110 -9782 20126 -9421
rect 20191 -9782 20216 -9421
rect 20110 -9799 20216 -9782
rect 26625 -9792 33073 -9388
rect 32669 -9861 33073 -9792
rect 26113 -10357 26150 -10331
rect 32660 -10732 33072 -10676
rect 26626 -11146 33073 -10732
rect 26635 -12182 33065 -11964
rect 26635 -12199 33006 -12182
rect 16200 -12616 16402 -12600
rect 16202 -12799 16402 -12616
rect 33400 -12418 33606 -12402
rect 33400 -12799 33598 -12418
rect 16180 -12997 16196 -12799
rect 33598 -12997 33614 -12799
rect 16202 -13000 16402 -12997
<< viali >>
rect 18320 -6069 18321 -5747
rect 18321 -6069 18455 -5747
rect 20392 -6067 20526 -5735
rect 20526 -6067 20528 -5735
rect 23740 -6548 23827 -4933
rect 24316 -4967 24386 -4932
rect 24316 -5200 24329 -4967
rect 24329 -5200 24372 -4967
rect 24372 -5200 24386 -4967
rect 26320 -4967 26390 -4898
rect 26320 -5166 26334 -4967
rect 26334 -5166 26377 -4967
rect 26377 -5166 26390 -4967
rect 24319 -6720 24329 -6221
rect 24329 -6720 24372 -6221
rect 24372 -6720 24387 -6221
rect 26321 -6724 26334 -6225
rect 26334 -6724 26377 -6225
rect 26377 -6724 26389 -6225
rect 16198 -8734 16200 -8094
rect 16200 -8734 16397 -8094
rect 16591 -8665 16594 -8116
rect 16594 -8665 16686 -8116
rect 16686 -8665 16687 -8116
rect 23824 -7749 23896 -7715
rect 23194 -8065 23235 -7834
rect 26076 -8099 26111 -7845
rect 22151 -8674 22154 -8125
rect 22154 -8674 22246 -8125
rect 22246 -8674 22247 -8125
rect 23196 -8845 23237 -8614
rect 26076 -8876 26111 -8622
rect 23492 -9007 23563 -8973
rect 18825 -9557 18890 -9426
rect 18825 -9787 18890 -9650
rect 20126 -9552 20191 -9421
rect 20126 -9782 20191 -9645
rect 23167 -9698 23204 -9305
rect 26112 -9700 26149 -9307
rect 23175 -10358 23212 -9965
rect 26113 -10331 26150 -9964
rect 23145 -12994 23259 -12880
rect 26061 -12980 26175 -12866
<< metal1 >>
rect 22521 -4257 26216 -4255
rect 22521 -4385 26158 -4257
rect 22521 -4496 22726 -4385
rect 26152 -4388 26158 -4385
rect 26289 -4388 26295 -4257
rect 22519 -4850 22726 -4496
rect 22382 -4854 22726 -4850
rect 23633 -4596 25934 -4500
rect 23633 -4700 25935 -4596
rect 18947 -5695 19923 -5692
rect 18266 -5747 18888 -5701
rect 18266 -6040 18320 -5747
rect 18268 -6069 18320 -6040
rect 18455 -5790 18888 -5747
rect 18947 -5755 19398 -5695
rect 19388 -5761 19398 -5755
rect 19483 -5755 19923 -5695
rect 19982 -5735 20599 -5701
rect 19483 -5761 19493 -5755
rect 19982 -5790 20392 -5735
rect 18455 -6067 20392 -5790
rect 20528 -6040 20599 -5735
rect 20528 -6067 20597 -6040
rect 18455 -6069 18558 -6067
rect 18314 -6081 18461 -6069
rect 20386 -6079 20534 -6067
rect 18888 -6768 18950 -6317
rect 19405 -6347 19467 -6300
rect 19378 -6505 19388 -6347
rect 19487 -6505 19497 -6347
rect 19404 -6599 19465 -6505
rect 19922 -6611 19984 -6314
rect 19922 -6734 21359 -6611
rect 21482 -6734 21488 -6611
rect 19343 -6768 19547 -6767
rect 19922 -6768 19984 -6734
rect 18888 -6830 19984 -6768
rect 19236 -6835 19547 -6830
rect 17618 -7029 17628 -6932
rect 17800 -7029 17832 -6932
rect 17628 -7733 17832 -7029
rect 19343 -7731 19547 -6835
rect 21539 -6838 21641 -4933
rect 22143 -6570 23155 -4854
rect 23633 -4933 23833 -4700
rect 24768 -4755 25935 -4700
rect 24323 -4815 24694 -4755
rect 24753 -4815 25959 -4755
rect 26018 -4815 26386 -4755
rect 24323 -4879 24383 -4815
rect 26326 -4878 26386 -4815
rect 26292 -4879 26412 -4878
rect 24299 -4880 26412 -4879
rect 23633 -6548 23740 -4933
rect 23827 -6548 23833 -4933
rect 24298 -4898 26412 -4880
rect 24298 -4932 26320 -4898
rect 24298 -5200 24316 -4932
rect 24386 -5166 26320 -4932
rect 26390 -5166 26412 -4898
rect 24386 -5200 26412 -5166
rect 24298 -5204 26412 -5200
rect 24298 -5206 24412 -5204
rect 26288 -5206 26412 -5204
rect 24298 -5208 24402 -5206
rect 24310 -5212 24392 -5208
rect 25775 -5976 26035 -5975
rect 26158 -5976 26288 -5970
rect 25775 -6106 26158 -5976
rect 24313 -6220 24393 -6209
rect 23633 -6671 23833 -6548
rect 23633 -6778 23756 -6671
rect 24308 -6720 24318 -6220
rect 24388 -6720 24590 -6220
rect 24313 -6732 24393 -6720
rect 21049 -7031 21059 -6925
rect 21267 -7031 21277 -6925
rect 21539 -6940 22240 -6838
rect 22367 -6901 22373 -6778
rect 22496 -6901 23756 -6778
rect 24816 -6935 24944 -6218
rect 21063 -7727 21267 -7031
rect 16192 -8094 16403 -8082
rect 16192 -8734 16198 -8094
rect 16397 -8201 16403 -8094
rect 16585 -8116 16693 -8104
rect 16585 -8122 16591 -8116
rect 16520 -8201 16591 -8122
rect 16397 -8601 16591 -8201
rect 16397 -8734 16403 -8601
rect 16192 -8746 16403 -8734
rect 16520 -8665 16591 -8601
rect 16687 -8132 16693 -8116
rect 22138 -8113 22240 -6940
rect 24812 -7121 24946 -6935
rect 22919 -7255 24946 -7121
rect 25146 -7183 25255 -6220
rect 22138 -8125 22253 -8113
rect 16687 -8665 17683 -8132
rect 16520 -8677 17683 -8665
rect 16520 -8784 16623 -8677
rect 16683 -8794 17683 -8677
rect 18486 -8195 20392 -8129
rect 22138 -8131 22151 -8125
rect 18486 -8644 18534 -8195
rect 18626 -8203 20392 -8195
rect 18626 -8644 20254 -8203
rect 18486 -8652 20254 -8644
rect 20346 -8652 20392 -8203
rect 18486 -8713 20392 -8652
rect 21183 -8674 22151 -8131
rect 22247 -8674 22253 -8125
rect 21183 -8686 22253 -8674
rect 18009 -8950 18178 -8742
rect 18608 -8753 20268 -8742
rect 18608 -8824 19789 -8753
rect 19783 -8853 19789 -8824
rect 19889 -8824 20268 -8753
rect 20654 -8746 20818 -8741
rect 19889 -8853 19895 -8824
rect 20654 -8846 20668 -8746
rect 20768 -8846 20818 -8746
rect 21183 -8793 22183 -8686
rect 20654 -8950 20818 -8846
rect 18009 -9097 20818 -8950
rect 18009 -9099 18178 -9097
rect 22919 -9175 23053 -7255
rect 25146 -7539 25255 -7292
rect 25454 -7374 25563 -6215
rect 25775 -7089 25893 -6106
rect 26158 -6112 26288 -6106
rect 26315 -6224 26395 -6213
rect 26132 -6723 26320 -6224
rect 26392 -6723 26402 -6224
rect 26132 -6724 26321 -6723
rect 26389 -6724 26402 -6723
rect 26315 -6736 26395 -6724
rect 25775 -7206 26356 -7089
rect 25775 -7207 26160 -7206
rect 25454 -7489 25563 -7483
rect 25146 -7624 25160 -7539
rect 25245 -7624 25815 -7539
rect 25146 -7626 25255 -7624
rect 25160 -7630 25245 -7626
rect 23812 -7715 23908 -7709
rect 23812 -7749 23824 -7715
rect 23896 -7749 23908 -7715
rect 23812 -7755 23908 -7749
rect 23255 -7799 23397 -7798
rect 23160 -7800 23397 -7799
rect 23140 -7834 23397 -7800
rect 23140 -8065 23194 -7834
rect 23235 -8065 23397 -7834
rect 23140 -8100 23397 -8065
rect 23493 -7845 23563 -7844
rect 23493 -8001 23729 -7845
rect 23140 -8469 23256 -8100
rect 23493 -8277 23563 -8001
rect 23659 -8278 23729 -8001
rect 23824 -8277 23896 -7755
rect 23991 -7809 24985 -7739
rect 23991 -8278 24061 -7809
rect 24156 -8001 24393 -7845
rect 24156 -8278 24226 -8001
rect 24323 -8278 24393 -8001
rect 24635 -8187 24684 -7880
rect 24626 -8239 24632 -8187
rect 24684 -8239 24690 -8187
rect 24635 -8246 24684 -8239
rect 24915 -8278 24985 -7809
rect 25081 -7809 25649 -7739
rect 25081 -8278 25151 -7809
rect 25247 -8001 25483 -7845
rect 25247 -8278 25317 -8001
rect 25413 -8278 25483 -8001
rect 25579 -8278 25649 -7809
rect 25730 -8273 25815 -7624
rect 25911 -7845 26147 -7832
rect 25911 -8099 26076 -7845
rect 26111 -8099 26147 -7845
rect 25911 -8100 26147 -8099
rect 25745 -8277 25815 -8273
rect 24618 -8422 24624 -8417
rect 23139 -8567 23256 -8469
rect 23139 -8588 23257 -8567
rect 23139 -8589 23397 -8588
rect 23138 -8614 23397 -8589
rect 23138 -8845 23196 -8614
rect 23237 -8845 23397 -8614
rect 23138 -8875 23397 -8845
rect 19402 -9247 19408 -9187
rect 19468 -9247 19474 -9187
rect 18819 -9421 18896 -9414
rect 18819 -9426 19145 -9421
rect 18819 -9557 18825 -9426
rect 18890 -9557 19145 -9426
rect 18819 -9558 19145 -9557
rect 18819 -9569 18896 -9558
rect 19408 -9561 19468 -9247
rect 19722 -9309 23053 -9175
rect 23139 -8877 23397 -8875
rect 23139 -8878 23297 -8877
rect 23139 -9297 23256 -8878
rect 23492 -8967 23563 -8501
rect 23659 -8906 23729 -8443
rect 23991 -8721 24061 -8443
rect 23825 -8877 24061 -8721
rect 24156 -8906 24226 -8443
rect 23480 -8973 23575 -8967
rect 23480 -9007 23492 -8973
rect 23563 -9007 23575 -8973
rect 23659 -8976 24226 -8906
rect 24323 -8908 24393 -8443
rect 24616 -8473 24624 -8422
rect 24680 -8422 24686 -8417
rect 24680 -8473 24691 -8422
rect 24616 -8830 24691 -8473
rect 24915 -8721 24985 -8436
rect 25081 -8721 25151 -8436
rect 24915 -8877 25151 -8721
rect 24915 -8878 24985 -8877
rect 25247 -8908 25317 -8436
rect 24323 -8978 25317 -8908
rect 25413 -8903 25483 -8447
rect 25579 -8721 25649 -8436
rect 26054 -8622 26147 -8100
rect 25579 -8877 25815 -8721
rect 25911 -8876 26076 -8622
rect 26111 -8876 26147 -8622
rect 25465 -8955 25483 -8903
rect 25911 -8910 26147 -8876
rect 25413 -8972 25483 -8955
rect 23480 -9013 23575 -9007
rect 26278 -9060 26356 -7206
rect 25658 -9131 26356 -9060
rect 25656 -9178 26356 -9131
rect 26925 -7285 32772 -4768
rect 26925 -8098 29439 -7285
rect 29528 -7600 30172 -7382
rect 29528 -7802 29809 -7600
rect 30011 -7802 30172 -7600
rect 29528 -8006 30172 -7802
rect 30255 -8098 32772 -7285
rect 26925 -8749 32772 -8098
rect 26925 -8799 29547 -8749
rect 29578 -8799 32772 -8749
rect 26925 -9000 32772 -8799
rect 25656 -9217 26023 -9178
rect 26925 -9200 29807 -9000
rect 30007 -9200 32772 -9000
rect 23139 -9305 23444 -9297
rect 18819 -9650 18915 -9638
rect 18794 -9787 18825 -9650
rect 18890 -9787 19624 -9650
rect 19722 -9747 19784 -9309
rect 20120 -9416 20197 -9409
rect 20120 -9421 20216 -9416
rect 20120 -9552 20126 -9421
rect 20191 -9552 20216 -9421
rect 20120 -9553 20216 -9552
rect 20120 -9564 20197 -9553
rect 18819 -9799 19162 -9787
rect 19251 -9794 19341 -9787
rect 18839 -9836 19162 -9799
rect 19662 -9809 19784 -9747
rect 19882 -9632 20103 -9631
rect 19882 -9645 20218 -9632
rect 19882 -9782 20126 -9645
rect 20191 -9653 20218 -9645
rect 20191 -9782 20219 -9653
rect 19882 -9797 20219 -9782
rect 23139 -9698 23167 -9305
rect 23204 -9310 23444 -9305
rect 23552 -9310 23671 -9297
rect 23204 -9698 23671 -9310
rect 23139 -9707 23671 -9698
rect 23139 -9708 23444 -9707
rect 18839 -9869 19254 -9836
rect 19662 -9841 19724 -9809
rect 19882 -9837 20218 -9797
rect 18843 -9891 19254 -9869
rect 19308 -9891 19725 -9841
rect 19778 -9891 20218 -9837
rect 23139 -9964 23256 -9708
rect 23552 -9725 23671 -9707
rect 23784 -9310 23903 -9299
rect 24019 -9310 24138 -9297
rect 23784 -9707 24138 -9310
rect 23784 -9725 23903 -9707
rect 24019 -9725 24138 -9707
rect 24254 -9313 24373 -9297
rect 24488 -9313 24607 -9298
rect 24254 -9710 24607 -9313
rect 24254 -9725 24373 -9710
rect 24488 -9725 24607 -9710
rect 24721 -9308 24840 -9298
rect 24955 -9308 25074 -9297
rect 24721 -9705 25074 -9308
rect 24721 -9725 24840 -9705
rect 24955 -9725 25074 -9705
rect 25190 -9311 25309 -9298
rect 25423 -9311 25542 -9298
rect 25190 -9708 25542 -9311
rect 25656 -9582 25776 -9217
rect 25891 -9261 26171 -9258
rect 25891 -9307 26181 -9261
rect 25891 -9394 26112 -9307
rect 25190 -9725 25309 -9708
rect 25423 -9725 25542 -9708
rect 25657 -9719 25776 -9582
rect 25897 -9700 26112 -9394
rect 26149 -9700 26181 -9307
rect 25897 -9705 26181 -9700
rect 23552 -9961 23671 -9945
rect 23784 -9961 23903 -9942
rect 23139 -9965 23433 -9964
rect 23139 -10358 23175 -9965
rect 23212 -10358 23433 -9965
rect 23139 -10359 23433 -10358
rect 23552 -10358 23903 -9961
rect 23139 -12880 23265 -10359
rect 23552 -10370 23671 -10358
rect 23784 -10372 23903 -10358
rect 24019 -9961 24138 -9942
rect 24254 -9961 24373 -9942
rect 24019 -10358 24373 -9961
rect 24019 -10370 24138 -10358
rect 24254 -10370 24373 -10358
rect 24488 -9961 24607 -9942
rect 24721 -9961 24840 -9942
rect 24488 -10358 24840 -9961
rect 24488 -10371 24607 -10358
rect 24721 -10371 24840 -10358
rect 24955 -9961 25074 -9942
rect 25190 -9961 25309 -9942
rect 24955 -10358 25309 -9961
rect 24955 -10370 25074 -10358
rect 25190 -10371 25309 -10358
rect 25423 -9963 25542 -9942
rect 25657 -9963 25776 -9945
rect 26088 -9963 26181 -9705
rect 25423 -10360 25776 -9963
rect 25896 -9964 26181 -9963
rect 25896 -10331 26113 -9964
rect 26150 -10331 26181 -9964
rect 25896 -10332 26181 -10331
rect 25423 -10371 25542 -10360
rect 25657 -10372 25776 -10360
rect 25889 -10512 26181 -10332
rect 23139 -12994 23145 -12880
rect 23259 -12994 23265 -12880
rect 26055 -12866 26181 -10512
rect 26925 -11902 32772 -9200
rect 26055 -12980 26061 -12866
rect 26175 -12980 26181 -12866
rect 26055 -12992 26181 -12980
rect 23139 -13006 23265 -12994
<< via1 >>
rect 26158 -4388 26289 -4257
rect 18320 -6069 18455 -5747
rect 19398 -5761 19483 -5695
rect 20392 -6067 20528 -5735
rect 19388 -6505 19487 -6347
rect 21359 -6734 21482 -6611
rect 17628 -7029 17800 -6932
rect 24316 -5200 24386 -4932
rect 26320 -5166 26390 -4898
rect 26158 -6106 26288 -5976
rect 24318 -6221 24388 -6220
rect 24318 -6720 24319 -6221
rect 24319 -6720 24387 -6221
rect 24387 -6720 24388 -6221
rect 21059 -7031 21267 -6925
rect 22373 -6901 22496 -6778
rect 18534 -8644 18626 -8195
rect 20254 -8652 20346 -8203
rect 19789 -8853 19889 -8753
rect 20668 -8846 20768 -8746
rect 25146 -7292 25255 -7183
rect 26320 -6225 26392 -6224
rect 26320 -6723 26321 -6225
rect 26321 -6723 26389 -6225
rect 26389 -6723 26392 -6225
rect 25454 -7483 25563 -7374
rect 25160 -7624 25245 -7539
rect 24632 -8239 24684 -8187
rect 19408 -9247 19468 -9187
rect 24624 -8473 24680 -8417
rect 25413 -8955 25465 -8903
rect 29809 -7802 30011 -7600
rect 29807 -9200 30007 -9000
<< metal2 >>
rect 26158 -4257 26289 -4251
rect 24316 -4932 24386 -4922
rect 24316 -5210 24386 -5200
rect 19398 -5695 19483 -5685
rect 18320 -5747 18455 -5737
rect 19398 -5771 19483 -5761
rect 20392 -5735 20528 -5725
rect 18320 -6079 18455 -6069
rect 19399 -6337 19473 -5771
rect 26158 -5976 26289 -4388
rect 26320 -4898 26390 -4888
rect 26320 -5176 26390 -5166
rect 20392 -6077 20528 -6067
rect 26152 -6106 26158 -5976
rect 26288 -6106 26294 -5976
rect 24318 -6220 24388 -6210
rect 19388 -6347 19487 -6337
rect 19388 -6515 19487 -6505
rect 17628 -6932 17800 -6922
rect 19399 -6950 19473 -6515
rect 21359 -6611 21482 -6605
rect 24318 -6730 24388 -6720
rect 26320 -6224 26392 -6214
rect 26320 -6733 26392 -6723
rect 21359 -6778 21482 -6734
rect 22373 -6778 22496 -6772
rect 21359 -6901 22373 -6778
rect 22373 -6907 22496 -6901
rect 21059 -6925 21267 -6915
rect 17800 -7024 21059 -6950
rect 17628 -7039 17800 -7029
rect 21059 -7041 21267 -7031
rect 25140 -7199 25146 -7183
rect 20668 -7292 25146 -7199
rect 25255 -7292 25261 -7183
rect 20668 -7299 25261 -7292
rect 18518 -8195 20374 -8155
rect 18518 -8644 18534 -8195
rect 18626 -8203 20374 -8195
rect 18626 -8644 20254 -8203
rect 18518 -8652 20254 -8644
rect 20346 -8652 20374 -8203
rect 18518 -8708 20374 -8652
rect 19364 -9187 19500 -8708
rect 20668 -8746 20768 -7299
rect 25448 -7397 25454 -7374
rect 19789 -8753 19889 -8747
rect 20668 -8852 20768 -8846
rect 22399 -7483 25454 -7397
rect 25563 -7397 25569 -7374
rect 26402 -7397 26604 -7394
rect 25563 -7483 26604 -7397
rect 22399 -7497 26604 -7483
rect 19789 -8901 19889 -8853
rect 22399 -8901 22499 -7497
rect 24621 -7624 25160 -7539
rect 25245 -7624 25251 -7539
rect 24621 -8187 24706 -7624
rect 24621 -8239 24632 -8187
rect 24684 -8239 24706 -8187
rect 24621 -8257 24706 -8239
rect 19789 -9001 22499 -8901
rect 24624 -8417 24680 -8411
rect 19364 -9247 19408 -9187
rect 19468 -9247 19500 -9187
rect 24624 -9006 24680 -8473
rect 25490 -8863 25538 -7497
rect 25566 -7502 25666 -7497
rect 26402 -7600 26604 -7497
rect 26402 -7802 29809 -7600
rect 30011 -7802 30017 -7600
rect 25413 -8903 25538 -8863
rect 25407 -8955 25413 -8903
rect 25465 -8953 25538 -8903
rect 25465 -8955 25471 -8953
rect 26400 -9000 26799 -8999
rect 26400 -9006 29807 -9000
rect 24624 -9196 29807 -9006
rect 26400 -9200 29807 -9196
rect 30007 -9200 30013 -9000
rect 19364 -9257 19500 -9247
<< via2 >>
rect 24316 -5200 24386 -4932
rect 18320 -6069 18455 -5747
rect 20392 -6067 20528 -5735
rect 26320 -5166 26390 -4898
rect 24318 -6720 24388 -6220
rect 26320 -6723 26392 -6224
<< metal3 >>
rect 20616 -4526 26396 -4525
rect 18315 -4703 26396 -4526
rect 18315 -4704 21394 -4703
rect 21818 -4704 26396 -4703
rect 18315 -4710 20636 -4704
rect 18315 -5742 18465 -4710
rect 20389 -5730 20526 -4710
rect 24312 -4927 24384 -4704
rect 26320 -4893 26392 -4704
rect 26310 -4898 26400 -4893
rect 24306 -4932 24396 -4927
rect 24306 -5200 24316 -4932
rect 24386 -5200 24396 -4932
rect 26310 -5166 26320 -4898
rect 26390 -5166 26400 -4898
rect 26310 -5171 26400 -5166
rect 24306 -5205 24396 -5200
rect 18310 -5747 18465 -5742
rect 18310 -6069 18320 -5747
rect 18455 -6069 18465 -5747
rect 18310 -6074 18465 -6069
rect 20382 -5735 20538 -5730
rect 20382 -6067 20392 -5735
rect 20528 -6067 20538 -5735
rect 20382 -6072 20538 -6067
rect 24312 -6215 24384 -5205
rect 24308 -6220 24398 -6215
rect 26320 -6219 26392 -5171
rect 24308 -6720 24318 -6220
rect 24388 -6720 24398 -6220
rect 24308 -6725 24398 -6720
rect 26310 -6224 26402 -6219
rect 26310 -6723 26320 -6224
rect 26392 -6723 26402 -6224
rect 24312 -6729 24384 -6725
rect 26310 -6728 26402 -6723
rect 26320 -6743 26392 -6728
use sky130_fd_pr__nfet_01v8_lvt_63HJ42  sky130_fd_pr__nfet_01v8_lvt_63HJ42_0
timestamp 1724943425
transform 1 0 19517 0 1 -9636
box -424 -257 424 257
use sky130_fd_pr__nfet_01v8_lvt_JQYUHL  sky130_fd_pr__nfet_01v8_lvt_JQYUHL_0
timestamp 1725314430
transform 1 0 19437 0 1 -7948
box -2603 -857 2603 857
use sky130_fd_pr__pfet_01v8_lvt_9BX3CZ  sky130_fd_pr__pfet_01v8_lvt_9BX3CZ_0
timestamp 1725314430
transform 1 0 19435 0 1 -6156
box -839 -498 839 464
use sky130_fd_pr__pfet_01v8_lvt_A7537V  sky130_fd_pr__pfet_01v8_lvt_A7537V_0
timestamp 1725314430
transform -1 0 22649 0 -1 -5723
box -1196 -973 1196 973
use sky130_fd_pr__res_xhigh_po_0p35_VRVSRL  sky130_fd_pr__res_xhigh_po_0p35_VRVSRL_0
timestamp 1724926688
transform -1 0 23860 0 -1 -8361
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p35_VUHUKX  sky130_fd_pr__res_xhigh_po_0p35_VUHUKX_0
timestamp 1725054279
transform -1 0 24654 0 -1 -8337
box -201 -672 201 672
use sky130_fd_pr__res_xhigh_po_0p35_Z5USRC  sky130_fd_pr__res_xhigh_po_0p35_Z5USRC_0
timestamp 1724926688
transform -1 0 25448 0 -1 -8361
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p69_5SXZXT  sky130_fd_pr__res_xhigh_po_0p69_5SXZXT_0
timestamp 1725054543
transform 1 0 24664 0 1 -9834
box -1522 -708 1522 708
use sky130_fd_pr__pfet_01v8_lvt_6GTY34  XM1
timestamp 1724939774
transform 1 0 25356 0 1 -5820
box -855 -1098 855 1064
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 5 1288
timestamp 1704896540
transform -1 0 33095 0 -1 -4445
box 0 0 1340 1340
<< labels >>
flabel metal3 20524 -4594 20654 -4534 0 FreeSans 320 0 0 0 VDD
port 1 nsew
rlabel metal2 23896 -7497 23996 -7397 1 MINUS
flabel metal1 22521 -4599 22724 -4401 0 FreeSans 160 0 0 0 Vbgr
port 2 nsew
flabel metal1 18986 -9776 19056 -9658 0 FreeSans 160 0 0 0 VSS
port 3 nsew
rlabel metal1 19409 -9364 19467 -9306 1 Sop
rlabel metal1 20061 -9272 20143 -9210 1 Gcm2
rlabel metal1 19928 -9309 20062 -9175 1 Gcm2
flabel metal1 22044 -8470 22115 -8196 0 FreeSans 160 0 0 0 VSS
port 3 nsew
flabel metal1 16413 -8587 16524 -8209 0 FreeSans 160 0 0 0 VSS
port 3 nsew
flabel metal1 19954 -9834 20043 -9662 0 FreeSans 160 0 0 0 VSS
port 3 nsew
rlabel nwell 19398 -6736 19475 -6628 1 Gcm1
flabel metal1 26278 -8396 26355 -8199 0 FreeSans 160 0 0 0 Vbgr
port 2 nsew
rlabel space 22487 -7298 22671 -7193 1 PLUS
flabel metal1 23163 -11573 23259 -11294 0 FreeSans 80 0 0 0 VSS
port 3 nsew
flabel metal1 26064 -11529 26162 -11132 0 FreeSans 80 0 0 0 VSS
port 3 nsew
flabel metal1 23148 -9136 23245 -9043 0 FreeSans 80 0 0 0 VSS
port 3 nsew
flabel metal1 22141 -7076 22232 -6950 0 FreeSans 80 0 0 0 VSS
port 3 nsew
<< end >>
