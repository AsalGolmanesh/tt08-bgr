magic
tech sky130A
magscale 1 2
timestamp 1724543890
<< pwell >>
rect -307 -3239 307 3239
<< psubdiff >>
rect -271 3169 -175 3203
rect 175 3169 271 3203
rect -271 3107 -237 3169
rect 237 3107 271 3169
rect -271 -3169 -237 -3107
rect 237 -3169 271 -3107
rect -271 -3203 -175 -3169
rect 175 -3203 271 -3169
<< psubdiffcont >>
rect -175 3169 175 3203
rect -271 -3107 -237 3107
rect 237 -3107 271 3107
rect -175 -3203 175 -3169
<< xpolycontact >>
rect -141 2641 141 3073
rect -141 -3073 141 -2641
<< xpolyres >>
rect -141 -2641 141 2641
<< locali >>
rect -271 3169 -175 3203
rect 175 3169 271 3203
rect -271 3107 -237 3169
rect 237 3107 271 3169
rect -271 -3169 -237 -3107
rect 237 -3169 271 -3107
rect -271 -3203 -175 -3169
rect 175 -3203 271 -3169
<< viali >>
rect -125 2658 125 3055
rect -125 -3055 125 -2658
<< metal1 >>
rect -131 3055 131 3067
rect -131 2658 -125 3055
rect 125 2658 131 3055
rect -131 2646 131 2658
rect -131 -2658 131 -2646
rect -131 -3055 -125 -2658
rect 125 -3055 131 -2658
rect -131 -3067 131 -3055
<< properties >>
string FIXED_BBOX -254 -3186 254 3186
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 26.57 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 37.954k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
