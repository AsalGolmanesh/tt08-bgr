magic
tech sky130A
magscale 1 2
timestamp 1725558127
<< viali >>
rect 6356 19182 7772 20010
<< metal1 >>
rect 6344 20010 7784 20016
rect 6344 19182 6356 20010
rect 7772 19182 7784 20010
rect 6344 19176 7784 19182
rect 18905 12278 20333 12421
rect 18866 9984 19042 10370
rect 19232 1860 19746 1908
rect 19176 1454 19186 1860
rect 19762 1823 19772 1860
rect 19762 1664 19846 1823
rect 20190 1664 20333 12278
rect 19762 1521 20333 1664
rect 19762 1454 19846 1521
rect 19187 1437 19846 1454
<< via1 >>
rect 6356 19182 7772 20010
rect 19186 1454 19762 1860
<< metal2 >>
rect 6356 20010 7772 20020
rect 6356 19172 7772 19182
rect 19186 1860 19762 1870
rect 19186 1444 19762 1454
<< via2 >>
rect 6356 19182 7772 20010
rect 19186 1454 19762 1860
<< metal3 >>
rect 6346 20010 7782 20015
rect 6346 19182 6356 20010
rect 7772 19182 7782 20010
rect 6346 19177 7782 19182
rect 5986 18010 8214 18054
rect 156 16646 176 18010
rect 578 17878 8214 18010
rect 578 16646 8266 17878
rect 156 16606 8266 16646
rect 5986 16580 8266 16606
rect 19176 1860 19772 1865
rect 19176 1454 19186 1860
rect 19762 1454 19772 1860
rect 19176 1449 19772 1454
<< via3 >>
rect 6356 19182 7772 20010
rect 176 16646 578 18010
rect 19186 1454 19762 1860
<< metal4 >>
rect 200 18011 600 44152
rect 800 44138 1200 44152
rect 6134 44138 6194 45152
rect 6686 44138 6746 45152
rect 7238 44138 7298 45152
rect 7790 44138 7850 45152
rect 8342 44138 8402 45152
rect 8894 44138 8954 45152
rect 9446 44138 9506 45152
rect 9998 44138 10058 45152
rect 10550 44138 10610 45152
rect 11102 44138 11162 45152
rect 11654 44138 11714 45152
rect 12206 44138 12266 45152
rect 12758 44138 12818 45152
rect 13310 44138 13370 45152
rect 13862 44138 13922 45152
rect 14414 44138 14474 45152
rect 14966 44138 15026 45152
rect 15518 44138 15578 45152
rect 16070 44138 16130 45152
rect 16622 44138 16682 45152
rect 17174 44138 17234 45152
rect 17726 44138 17786 45152
rect 18278 44138 18338 45152
rect 18830 44138 18890 45152
rect 19382 44936 19442 45152
rect 19934 44936 19994 45152
rect 20486 44936 20546 45152
rect 21038 44936 21098 45152
rect 21590 44936 21650 45152
rect 22142 44936 22202 45152
rect 22694 44936 22754 45152
rect 23246 44936 23306 45152
rect 23798 44936 23858 45152
rect 24350 44936 24410 45152
rect 24902 44936 24962 45152
rect 25454 44936 25514 45152
rect 26006 44936 26066 45152
rect 26558 44936 26618 45152
rect 27110 44936 27170 45152
rect 27662 44936 27722 45152
rect 28214 44936 28274 45152
rect 28766 44936 28826 45152
rect 29318 44916 29378 45152
rect 800 44134 19296 44138
rect 800 42930 29814 44134
rect 800 20010 1200 42930
rect 6355 20010 7773 20011
rect 794 19182 6356 20010
rect 7772 19182 8426 20010
rect 794 19028 8426 19182
rect 175 18010 600 18011
rect 175 16646 176 18010
rect 578 16646 600 18010
rect 175 16645 600 16646
rect 200 1000 600 16645
rect 800 5188 1200 19028
rect 800 2702 1196 5188
rect 800 1000 1200 2702
rect 19185 1860 19763 1861
rect 19185 1650 19186 1860
rect 18770 1470 19186 1650
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 1470
rect 19185 1454 19186 1470
rect 19762 1454 19763 1860
rect 19185 1453 19763 1454
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use core_prel  core_prel_0
timestamp 1725529118
transform 1 0 -2050 0 1 23047
box 6004 -19007 24007 -2979
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel space 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 800 5188 1200 44152 0 FreeSans 800 0 0 0 VGND
port 54 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
