magic
tech sky130A
magscale 1 2
timestamp 1724543890
<< error_s >>
rect -41 48 -6 82
rect -40 29 -6 48
rect -370 -2227 -355 -949
rect -336 -2227 -302 -895
rect -336 -2261 -321 -2227
rect -21 -2280 -6 29
rect 13 -5 48 29
rect 13 -2280 47 -5
rect 13 -2314 28 -2280
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__pfet_01v8_lvt_SX4MVH  XM1
timestamp 1724543890
transform 1 0 5380 0 1 1767
box -246 -2219 246 2219
use sky130_fd_pr__pfet_01v8_lvt_SX4MVH  XM2
timestamp 1724543890
transform 1 0 6470 0 1 1767
box -246 -2219 246 2219
use sky130_fd_pr__pfet_01v8_lvt_SX4MVH  XM3
timestamp 1724543890
transform 1 0 7526 0 1 1861
box -246 -2219 246 2219
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1704896540
transform 1 0 578 0 1 2768
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2
array 0 2 1288 0 10 1288
timestamp 1704896540
transform 1 0 -1968 0 1 5000
box 0 0 1340 1340
use sky130_fd_pr__res_xhigh_po_1p41_NPWLJD  XR1
timestamp 1724543890
transform 1 0 3529 0 1 2421
box -307 -3239 307 3239
use sky130_fd_pr__res_xhigh_po_0p35_HU4QAP  XR2
timestamp 1724543890
transform 1 0 -171 0 1 -1099
box -201 -1217 201 1217
use sky130_fd_pr__res_xhigh_po_0p35_HU4QAP  XR3
timestamp 1724543890
transform 1 0 178 0 1 -1152
box -201 -1217 201 1217
use sky130_fd_pr__res_xhigh_po_0p35_YK563K  XR19
timestamp 1724543890
transform 1 0 -520 0 1 -1588
box -201 -675 201 675
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 MINUS
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 PLUS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vbgr
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vp
<< end >>
