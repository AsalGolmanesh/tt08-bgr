magic
tech sky130A
magscale 1 2
timestamp 1725036214
<< nwell >>
rect 24100 -4757 24530 -4756
rect 18919 -7120 19291 -5355
rect 20451 -7120 20883 -5358
rect 24100 -6921 24702 -4757
rect 26205 -6494 26499 -4753
rect 26188 -6918 26499 -6494
rect 20706 -7121 20883 -7120
<< pwell >>
rect 23884 -7845 23954 -7746
rect 24974 -7845 25044 -7739
rect 25638 -7873 25708 -7823
rect 23071 -8122 23136 -8091
rect 23140 -8878 23190 -8621
rect 24216 -8978 24286 -8877
rect 25306 -8978 25376 -8877
rect 23060 -9808 23127 -9581
rect 23105 -10359 23326 -9964
<< nbase >>
rect 29575 -9292 29614 -9291
<< pdiff >>
rect 29575 -9292 29614 -9291
<< psubdiff >>
rect 16171 -3802 16195 -3600
rect 33602 -3802 33626 -3600
rect 16200 -4004 16402 -3980
rect 33402 -4202 33606 -4178
rect 16900 -7475 17099 -7399
rect 16900 -8923 16943 -7475
rect 17049 -8923 17099 -7475
rect 16900 -9002 17099 -8923
rect 22599 -7469 22798 -7393
rect 22599 -8917 22642 -7469
rect 22748 -8917 22798 -7469
rect 22599 -8996 22798 -8917
rect 19198 -9426 19404 -9399
rect 19198 -9787 19258 -9426
rect 19323 -9787 19404 -9426
rect 19198 -9800 19404 -9787
rect 20501 -9421 20707 -9394
rect 20501 -9782 20561 -9421
rect 20626 -9782 20707 -9421
rect 20501 -9795 20707 -9782
rect 33402 -12426 33606 -12402
rect 16200 -12624 16402 -12600
rect 16172 -12997 16196 -12799
rect 33598 -12997 33622 -12799
<< nsubdiff >>
rect 24300 -4967 24403 -4901
rect 19067 -5457 19216 -5403
rect 19067 -6902 19097 -5457
rect 19184 -6902 19216 -5457
rect 19067 -7004 19216 -6902
rect 20500 -5457 20649 -5398
rect 20500 -6902 20528 -5457
rect 20615 -6902 20649 -5457
rect 24300 -6747 24329 -4967
rect 24372 -6747 24403 -4967
rect 24300 -6802 24403 -6747
rect 26305 -4967 26408 -4901
rect 26305 -6747 26334 -4967
rect 26377 -6747 26408 -4967
rect 26305 -6802 26408 -6747
rect 20500 -6999 20649 -6902
<< psubdiffcont >>
rect 16195 -3802 33602 -3600
rect 16200 -12600 16402 -4004
rect 16943 -8923 17049 -7475
rect 22642 -8917 22748 -7469
rect 19258 -9787 19323 -9426
rect 20561 -9782 20626 -9421
rect 33402 -12402 33606 -4202
rect 16196 -12997 33598 -12799
<< nsubdiffcont >>
rect 19097 -6902 19184 -5457
rect 20528 -6902 20615 -5457
rect 24329 -6747 24372 -4967
rect 26334 -6747 26377 -4967
<< locali >>
rect 16179 -3802 16195 -3600
rect 33602 -3802 33618 -3600
rect 16202 -3988 16402 -3802
rect 16200 -4004 16402 -3988
rect 33400 -4100 33602 -3802
rect 33400 -4174 33606 -4100
rect 33402 -4202 33606 -4174
rect 26630 -4488 33006 -4471
rect 26630 -4707 33070 -4488
rect 19084 -5457 19197 -5429
rect 19084 -5467 19097 -5457
rect 19184 -5467 19197 -5457
rect 20518 -5457 20631 -5433
rect 19084 -5969 19086 -5467
rect 20518 -5472 20528 -5457
rect 20615 -5472 20631 -5457
rect 19084 -6902 19097 -5969
rect 19184 -6902 19197 -5969
rect 19084 -6954 19197 -6902
rect 20518 -5974 20521 -5472
rect 20518 -6902 20528 -5974
rect 20615 -6902 20631 -5974
rect 24317 -6747 24329 -5200
rect 24372 -6747 24384 -5200
rect 24317 -6784 24384 -6747
rect 26322 -6747 26334 -5200
rect 26377 -6747 26389 -5200
rect 26631 -5996 33071 -5523
rect 26322 -6784 26389 -6747
rect 20518 -6958 20631 -6902
rect 26630 -7284 33073 -6813
rect 16929 -7475 17070 -7444
rect 16929 -8923 16943 -7475
rect 17049 -8923 17070 -7475
rect 16929 -8926 16960 -8923
rect 17029 -8926 17070 -8923
rect 16929 -8973 17070 -8926
rect 22628 -7469 22769 -7438
rect 22628 -8917 22642 -7469
rect 22748 -8917 22769 -7469
rect 26627 -8572 33072 -8099
rect 22628 -8967 22769 -8917
rect 29575 -9292 29614 -9291
rect 19242 -9426 19348 -9401
rect 19242 -9787 19258 -9426
rect 19323 -9787 19348 -9426
rect 19242 -9804 19348 -9787
rect 20545 -9421 20651 -9396
rect 20545 -9651 20561 -9421
rect 20545 -9782 20560 -9651
rect 20626 -9782 20651 -9421
rect 20545 -9795 20651 -9782
rect 26625 -9792 33073 -9388
rect 32669 -9861 33073 -9792
rect 26006 -10357 26043 -10331
rect 32660 -10732 33072 -10676
rect 26626 -11146 33073 -10732
rect 26635 -12182 33065 -11964
rect 26635 -12199 33006 -12182
rect 16200 -12616 16402 -12600
rect 16202 -12799 16402 -12616
rect 33400 -12418 33606 -12402
rect 33400 -12799 33598 -12418
rect 16180 -12997 16196 -12799
rect 33598 -12997 33614 -12799
rect 16202 -13000 16402 -12997
<< viali >>
rect 19086 -5969 19097 -5467
rect 19097 -5969 19184 -5467
rect 19184 -5969 19198 -5467
rect 20521 -5974 20528 -5472
rect 20528 -5974 20615 -5472
rect 20615 -5974 20633 -5472
rect 21440 -6577 21498 -4880
rect 24316 -4967 24386 -4932
rect 24316 -5200 24329 -4967
rect 24329 -5200 24372 -4967
rect 24372 -5200 24386 -4967
rect 26320 -4967 26390 -4898
rect 26320 -5166 26334 -4967
rect 26334 -5166 26377 -4967
rect 26377 -5166 26390 -4967
rect 16204 -7774 16402 -7506
rect 16402 -7774 16472 -7506
rect 16960 -8923 17029 -7506
rect 16960 -8926 17029 -8923
rect 22655 -8909 22724 -7489
rect 23717 -7749 23789 -7715
rect 23087 -8065 23128 -7834
rect 25969 -8099 26004 -7845
rect 23075 -8324 23126 -8107
rect 23089 -8845 23130 -8614
rect 25969 -8876 26004 -8622
rect 23385 -9007 23456 -8973
rect 19258 -9557 19323 -9426
rect 19258 -9787 19323 -9650
rect 20560 -9782 20561 -9651
rect 20561 -9782 20626 -9651
rect 23060 -9698 23097 -9305
rect 26005 -9700 26042 -9307
rect 23068 -10358 23105 -9965
rect 26006 -10331 26043 -9964
rect 23038 -12985 23152 -12871
rect 25954 -12987 26068 -12873
<< metal1 >>
rect 22344 -4257 26216 -4255
rect 22344 -4385 26158 -4257
rect 22344 -4388 22550 -4385
rect 26152 -4388 26158 -4385
rect 26289 -4388 26295 -4257
rect 22344 -4496 22549 -4388
rect 22343 -4637 22549 -4496
rect 24068 -4631 24074 -4502
rect 24203 -4503 24216 -4502
rect 24203 -4631 24231 -4503
rect 21407 -4880 21610 -4745
rect 19112 -5416 19584 -5360
rect 19641 -5361 20101 -5357
rect 19641 -5410 19700 -5361
rect 19654 -5411 19700 -5410
rect 19112 -5455 19168 -5416
rect 19690 -5418 19700 -5411
rect 19800 -5410 20101 -5361
rect 19800 -5418 19810 -5410
rect 20155 -5417 20593 -5370
rect 19080 -5467 19204 -5455
rect 20546 -5460 20593 -5417
rect 19080 -5969 19086 -5467
rect 19198 -5470 19204 -5467
rect 20515 -5470 20639 -5460
rect 19198 -5472 20639 -5470
rect 19198 -5969 20521 -5472
rect 19080 -5972 20521 -5969
rect 19080 -5981 19204 -5972
rect 20515 -5974 20521 -5972
rect 20633 -5974 20639 -5472
rect 20515 -5986 20639 -5974
rect 19590 -6589 19636 -6533
rect 19588 -6595 19690 -6589
rect 19588 -6703 19690 -6697
rect 19590 -7083 19636 -6703
rect 18990 -7129 19636 -7083
rect 20106 -7081 20152 -6536
rect 21407 -6577 21440 -4880
rect 21498 -6577 21610 -4880
rect 22343 -4896 22551 -4637
rect 24201 -4670 24231 -4631
rect 24201 -4700 25934 -4670
rect 24769 -4755 24836 -4700
rect 24928 -4755 24995 -4700
rect 25083 -4755 25150 -4700
rect 25239 -4755 25306 -4700
rect 25403 -4755 25470 -4700
rect 25558 -4755 25625 -4700
rect 25713 -4755 25780 -4700
rect 25867 -4755 25934 -4700
rect 24323 -4815 24694 -4755
rect 24753 -4815 25959 -4755
rect 26018 -4815 26386 -4755
rect 24323 -4879 24383 -4815
rect 26326 -4878 26386 -4815
rect 26292 -4879 26412 -4878
rect 24299 -4880 26412 -4879
rect 21956 -6574 22957 -4896
rect 24298 -4898 26412 -4880
rect 24298 -4932 26320 -4898
rect 21407 -6691 21610 -6577
rect 21551 -7070 21606 -6691
rect 23614 -6775 23668 -4961
rect 24298 -5200 24316 -4932
rect 24386 -5166 26320 -4932
rect 26390 -5166 26412 -4898
rect 24386 -5200 26412 -5166
rect 24298 -5204 26412 -5200
rect 24298 -5206 24412 -5204
rect 26288 -5206 26412 -5204
rect 24298 -5208 24402 -5206
rect 24310 -5212 24392 -5208
rect 26158 -5976 26288 -5970
rect 25808 -6106 26158 -5976
rect 22666 -6829 23668 -6775
rect 22119 -7040 22468 -6913
rect 22595 -7040 22601 -6913
rect 22119 -7060 22238 -7040
rect 21784 -7070 22238 -7060
rect 20916 -7080 22238 -7070
rect 20705 -7081 22238 -7080
rect 20106 -7127 22238 -7081
rect 16954 -7500 17035 -7494
rect 16192 -7506 17309 -7500
rect 16192 -7774 16204 -7506
rect 16472 -7774 16960 -7506
rect 16192 -7780 16960 -7774
rect 16946 -7801 16960 -7780
rect 16954 -8926 16960 -7801
rect 17029 -7801 17309 -7506
rect 17029 -8926 17035 -7801
rect 18990 -7867 19036 -7129
rect 20705 -7155 22238 -7127
rect 20706 -7851 20752 -7155
rect 20916 -7163 22238 -7155
rect 21784 -7171 22238 -7163
rect 22666 -7469 22720 -6829
rect 24859 -7158 24905 -6219
rect 25176 -7098 25224 -6218
rect 25176 -7146 25379 -7098
rect 22830 -7277 24905 -7158
rect 25331 -7200 25379 -7146
rect 25492 -7200 25537 -6219
rect 25808 -7000 25857 -6106
rect 26158 -6112 26288 -6106
rect 25804 -7156 25861 -7000
rect 25331 -7203 25387 -7200
rect 22666 -7477 22724 -7469
rect 22649 -7489 22730 -7477
rect 22649 -7502 22655 -7489
rect 22403 -7803 22655 -7502
rect 20706 -7853 20712 -7851
rect 20746 -7853 20752 -7851
rect 20706 -7865 20752 -7853
rect 22649 -8099 22655 -7803
rect 22636 -8340 22655 -8099
rect 19829 -8446 19839 -8445
rect 18126 -8701 19839 -8446
rect 19905 -8446 19915 -8445
rect 19905 -8447 21608 -8446
rect 19905 -8701 21609 -8447
rect 16954 -8938 17035 -8926
rect 16964 -8988 17028 -8938
rect 21584 -8943 21609 -8701
rect 22649 -8909 22655 -8340
rect 22724 -8099 22730 -7489
rect 22830 -7569 22964 -7277
rect 25289 -7301 25299 -7203
rect 25377 -7301 25387 -7203
rect 25492 -7245 25694 -7200
rect 22823 -7703 22829 -7569
rect 22963 -7703 22969 -7569
rect 25331 -7572 25379 -7301
rect 25649 -7391 25694 -7245
rect 25799 -7299 26290 -7156
rect 26925 -7285 32772 -4768
rect 25594 -7397 25694 -7391
rect 25594 -7503 25694 -7497
rect 25329 -7578 25381 -7572
rect 25649 -7592 25694 -7503
rect 25329 -7636 25381 -7630
rect 23705 -7715 23801 -7709
rect 23705 -7749 23717 -7715
rect 23789 -7749 23801 -7715
rect 23705 -7755 23801 -7749
rect 23053 -7834 23148 -7799
rect 23053 -8065 23087 -7834
rect 23128 -7845 23148 -7834
rect 23386 -7845 23456 -7844
rect 23128 -8065 23290 -7845
rect 23053 -8099 23290 -8065
rect 22724 -8100 23290 -8099
rect 23386 -8001 23622 -7845
rect 22724 -8107 23149 -8100
rect 22724 -8324 23075 -8107
rect 23126 -8324 23149 -8107
rect 23386 -8277 23456 -8001
rect 22724 -8340 23149 -8324
rect 22724 -8909 22730 -8340
rect 22649 -8921 22730 -8909
rect 23053 -8567 23149 -8340
rect 23053 -8614 23150 -8567
rect 23053 -8845 23089 -8614
rect 23130 -8621 23150 -8614
rect 23130 -8845 23290 -8621
rect 23053 -8877 23290 -8845
rect 23053 -8878 23190 -8877
rect 16964 -9052 18112 -8988
rect 19694 -8992 19704 -8960
rect 18181 -9048 19704 -8992
rect 19800 -9048 19810 -8960
rect 19990 -8992 20000 -8960
rect 19931 -9048 20000 -8992
rect 20100 -8992 20110 -8960
rect 20100 -9048 21555 -8992
rect 22667 -8994 22724 -8921
rect 21611 -9051 22724 -8994
rect 19835 -9247 19841 -9187
rect 19901 -9247 19907 -9187
rect 21418 -9211 22829 -9175
rect 19252 -9421 19329 -9414
rect 19252 -9426 19578 -9421
rect 19252 -9557 19258 -9426
rect 19323 -9557 19578 -9426
rect 19252 -9558 19578 -9557
rect 19252 -9569 19329 -9558
rect 19841 -9561 19901 -9247
rect 20155 -9273 22829 -9211
rect 19252 -9650 19348 -9638
rect 19227 -9787 19258 -9650
rect 19323 -9787 20057 -9650
rect 20155 -9747 20217 -9273
rect 21418 -9309 22829 -9273
rect 22963 -9309 22969 -9175
rect 23053 -9300 23149 -8878
rect 23385 -8967 23456 -8445
rect 23552 -8906 23622 -8001
rect 23717 -8277 23789 -7755
rect 23884 -7809 24878 -7739
rect 23884 -8721 23954 -7809
rect 23718 -8877 23954 -8721
rect 24049 -8001 24286 -7845
rect 24049 -8906 24119 -8001
rect 23373 -8973 23468 -8967
rect 23373 -9007 23385 -8973
rect 23456 -9007 23468 -8973
rect 23552 -8976 24119 -8906
rect 24216 -8908 24286 -8001
rect 24509 -8830 24519 -8422
rect 24574 -8830 24584 -8422
rect 24808 -8721 24878 -7809
rect 24974 -7809 25542 -7739
rect 24974 -8721 25044 -7809
rect 24808 -8877 25044 -8721
rect 25140 -8001 25376 -7845
rect 24808 -8878 24878 -8877
rect 25140 -8908 25210 -8001
rect 24216 -8978 25210 -8908
rect 25306 -8903 25376 -8001
rect 25472 -8721 25542 -7809
rect 25638 -8277 25708 -7592
rect 25963 -7845 26010 -7833
rect 25804 -8099 25969 -7845
rect 26004 -8099 26010 -7845
rect 26170 -8011 26289 -7299
rect 25804 -8100 26010 -8099
rect 25963 -8111 26010 -8100
rect 25963 -8622 26010 -8610
rect 25472 -8877 25708 -8721
rect 25804 -8876 25969 -8622
rect 26004 -8876 26010 -8622
rect 25804 -8877 26010 -8876
rect 25963 -8888 26010 -8877
rect 25358 -8955 25376 -8903
rect 25306 -8978 25376 -8955
rect 23373 -9013 23468 -9007
rect 26171 -9078 26289 -8011
rect 26170 -9098 26289 -9078
rect 25549 -9217 26289 -9098
rect 26925 -8098 29439 -7285
rect 29528 -8006 29538 -7382
rect 30162 -8006 30172 -7382
rect 30255 -8098 32772 -7285
rect 26925 -8654 32772 -8098
rect 26925 -8749 29588 -8654
rect 26925 -8799 29547 -8749
rect 29578 -8799 29588 -8749
rect 23053 -9305 23150 -9300
rect 20554 -9651 20632 -9639
rect 19252 -9793 19348 -9787
rect 19252 -9799 19341 -9793
rect 19684 -9794 19774 -9787
rect 19276 -9836 19341 -9799
rect 20095 -9809 20217 -9747
rect 20322 -9782 20560 -9651
rect 20626 -9782 20652 -9651
rect 20322 -9788 20652 -9782
rect 23053 -9698 23060 -9305
rect 23097 -9533 23150 -9305
rect 23200 -9310 23262 -9300
rect 23445 -9310 23564 -9297
rect 23200 -9533 23564 -9310
rect 23097 -9698 23149 -9533
rect 20554 -9794 20632 -9788
rect 19276 -9899 19687 -9836
rect 20095 -9841 20157 -9809
rect 20561 -9837 20626 -9794
rect 19741 -9899 20158 -9841
rect 20215 -9900 20626 -9837
rect 23053 -9954 23149 -9698
rect 23216 -9707 23564 -9533
rect 23445 -9725 23564 -9707
rect 23677 -9310 23796 -9299
rect 23912 -9310 24031 -9297
rect 23677 -9707 24031 -9310
rect 23032 -9964 23158 -9954
rect 23445 -9961 23564 -9945
rect 23677 -9961 23796 -9707
rect 23032 -9965 23326 -9964
rect 23032 -10358 23068 -9965
rect 23105 -10358 23326 -9965
rect 23032 -10359 23326 -10358
rect 23445 -10358 23796 -9961
rect 23032 -12871 23158 -10359
rect 23445 -10370 23564 -10358
rect 23677 -10372 23796 -10358
rect 23912 -9961 24031 -9707
rect 24147 -9313 24266 -9297
rect 24381 -9313 24500 -9298
rect 24147 -9710 24500 -9313
rect 24147 -9961 24266 -9710
rect 23912 -10358 24266 -9961
rect 23912 -10370 24031 -10358
rect 24147 -10370 24266 -10358
rect 24381 -9961 24500 -9710
rect 24614 -9308 24733 -9298
rect 24848 -9308 24967 -9297
rect 24614 -9705 24967 -9308
rect 24614 -9961 24733 -9705
rect 24381 -10358 24733 -9961
rect 24381 -10371 24500 -10358
rect 24614 -10371 24733 -10358
rect 24848 -9961 24967 -9705
rect 25083 -9311 25202 -9298
rect 25316 -9311 25435 -9298
rect 25083 -9708 25435 -9311
rect 25549 -9299 25668 -9217
rect 25549 -9582 25669 -9299
rect 25999 -9307 26048 -9295
rect 25999 -9310 26005 -9307
rect 25083 -9961 25202 -9708
rect 24848 -10358 25202 -9961
rect 24848 -10370 24967 -10358
rect 25083 -10371 25202 -10358
rect 25316 -9963 25435 -9708
rect 25550 -9719 25669 -9582
rect 25790 -9700 26005 -9310
rect 26042 -9700 26048 -9307
rect 25790 -9705 26048 -9700
rect 25999 -9712 26048 -9705
rect 26925 -9298 29588 -8799
rect 30186 -9298 32772 -8654
rect 25550 -9963 25669 -9945
rect 26002 -9952 26074 -9948
rect 26000 -9963 26074 -9952
rect 25316 -10360 25669 -9963
rect 25789 -9964 26074 -9963
rect 25789 -10331 26006 -9964
rect 26043 -10331 26074 -9964
rect 25789 -10357 26074 -10331
rect 25789 -10358 25918 -10357
rect 25316 -10371 25435 -10360
rect 25550 -10372 25669 -10360
rect 23032 -12985 23038 -12871
rect 23152 -12985 23158 -12871
rect 23032 -12997 23158 -12985
rect 25948 -12873 26074 -10357
rect 26925 -11902 32772 -9298
rect 25948 -12987 25954 -12873
rect 26068 -12987 26074 -12873
rect 25948 -12999 26074 -12987
<< via1 >>
rect 26158 -4388 26289 -4257
rect 24074 -4631 24203 -4502
rect 19700 -5418 19800 -5361
rect 19090 -5918 19182 -5480
rect 20526 -5916 20618 -5478
rect 19588 -6697 19690 -6595
rect 24316 -5200 24386 -4932
rect 26320 -5166 26390 -4898
rect 26158 -6106 26288 -5976
rect 22468 -7040 22595 -6913
rect 19839 -8701 19905 -8445
rect 25299 -7301 25377 -7203
rect 22829 -7703 22963 -7569
rect 25594 -7497 25694 -7397
rect 25329 -7630 25381 -7578
rect 19704 -9048 19800 -8960
rect 20000 -9048 20100 -8960
rect 19841 -9247 19901 -9187
rect 22829 -9309 22963 -9175
rect 24519 -8830 24574 -8422
rect 25306 -8955 25358 -8903
rect 29538 -8006 30162 -7382
rect 29588 -9298 30186 -8654
<< metal2 >>
rect 26158 -4257 26289 -4251
rect 24074 -4502 24203 -4496
rect 19700 -5361 19800 -5351
rect 19700 -5438 19800 -5418
rect 19090 -5480 19182 -5470
rect 19090 -5928 19182 -5918
rect 19700 -6595 19802 -5438
rect 20526 -5478 20618 -5468
rect 20526 -5926 20618 -5916
rect 19582 -6697 19588 -6595
rect 19690 -6697 19802 -6595
rect 22468 -6910 22595 -6907
rect 24074 -6910 24203 -4631
rect 24316 -4932 24386 -4922
rect 24316 -5210 24386 -5200
rect 26158 -5976 26289 -4388
rect 26320 -4898 26390 -4888
rect 26320 -5176 26390 -5166
rect 26152 -6106 26158 -5976
rect 26288 -6106 26294 -5976
rect 22468 -6913 24203 -6910
rect 22595 -7040 24203 -6913
rect 22468 -7046 22595 -7040
rect 25299 -7199 25380 -7193
rect 19704 -7203 25380 -7199
rect 19704 -7299 25299 -7203
rect 19704 -8960 19804 -7299
rect 25377 -7299 25380 -7203
rect 25299 -7311 25377 -7301
rect 29538 -7382 30162 -7372
rect 20001 -7497 25594 -7397
rect 25694 -7497 25700 -7397
rect 26286 -7467 29538 -7382
rect 19839 -8445 19905 -8435
rect 19839 -8711 19905 -8701
rect 19840 -8950 19902 -8711
rect 20001 -8950 20101 -7497
rect 19800 -9040 19804 -8960
rect 19704 -9058 19800 -9048
rect 19841 -9187 19901 -8950
rect 20000 -8960 20101 -8950
rect 20100 -9043 20101 -8960
rect 22829 -7569 22963 -7563
rect 26287 -7578 29538 -7467
rect 25323 -7630 25329 -7578
rect 25381 -7630 29538 -7578
rect 25400 -7634 29538 -7630
rect 20000 -9058 20100 -9048
rect 19841 -9253 19901 -9247
rect 22829 -9175 22963 -7703
rect 24512 -8422 24582 -8411
rect 24512 -8830 24519 -8422
rect 24574 -8830 24582 -8422
rect 24512 -9033 24582 -8830
rect 25300 -8955 25306 -8903
rect 25358 -8905 25364 -8903
rect 25402 -8905 25450 -7634
rect 26333 -7922 29538 -7634
rect 26595 -8006 29538 -7922
rect 29538 -8016 30162 -8006
rect 29588 -8654 30186 -8644
rect 29503 -8667 29588 -8665
rect 26594 -8718 29588 -8667
rect 26595 -8749 29588 -8718
rect 25358 -8953 25450 -8905
rect 25358 -8955 25364 -8953
rect 26328 -9033 29588 -8749
rect 24512 -9103 29588 -9033
rect 26187 -9206 29588 -9103
rect 26188 -9291 29588 -9206
rect 30186 -9289 30191 -8665
rect 29588 -9308 30186 -9298
rect 22829 -9315 22963 -9309
<< via2 >>
rect 19090 -5918 19182 -5480
rect 20526 -5916 20618 -5478
rect 24316 -5200 24386 -4932
rect 26320 -5166 26390 -4898
<< metal3 >>
rect 19104 -4598 26392 -4526
rect 19104 -5475 19176 -4598
rect 20532 -5473 20604 -4598
rect 24312 -4927 24384 -4598
rect 26320 -4893 26392 -4598
rect 26310 -4898 26400 -4893
rect 24306 -4932 24396 -4927
rect 24306 -5200 24316 -4932
rect 24386 -5200 24396 -4932
rect 26310 -5166 26320 -4898
rect 26390 -5166 26400 -4898
rect 26310 -5171 26400 -5166
rect 24306 -5205 24396 -5200
rect 19080 -5480 19192 -5475
rect 19080 -5918 19090 -5480
rect 19182 -5918 19192 -5480
rect 19080 -5923 19192 -5918
rect 20516 -5478 20628 -5473
rect 20516 -5916 20526 -5478
rect 20618 -5916 20628 -5478
rect 20516 -5921 20628 -5916
rect 20532 -5966 20604 -5921
use sky130_fd_pr__nfet_01v8_lvt_63HJ42  sky130_fd_pr__nfet_01v8_lvt_63HJ42_0
timestamp 1724943425
transform 1 0 19950 0 1 -9636
box -424 -257 424 257
use sky130_fd_pr__nfet_01v8_lvt_JUYCGL  sky130_fd_pr__nfet_01v8_lvt_JUYCGL_0
timestamp 1724941373
transform 1 0 19868 0 1 -8191
box -2603 -857 2603 857
use sky130_fd_pr__pfet_01v8_lvt_W4537V  sky130_fd_pr__pfet_01v8_lvt_W4537V_0
timestamp 1725004556
transform -1 0 22610 0 -1 -5723
box -1196 -973 1196 973
use sky130_fd_pr__pfet_01v8_W45NJQ  sky130_fd_pr__pfet_01v8_W45NJQ_0
timestamp 1724940898
transform 1 0 19871 0 1 -6222
box -581 -898 581 864
use sky130_fd_pr__res_xhigh_po_0p35_PZL4NP  sky130_fd_pr__res_xhigh_po_0p35_PZL4NP_0
timestamp 1724945390
transform -1 0 24547 0 -1 -8337
box -201 -672 201 672
use sky130_fd_pr__res_xhigh_po_0p35_VRVSRL  sky130_fd_pr__res_xhigh_po_0p35_VRVSRL_0
timestamp 1724926688
transform -1 0 23753 0 -1 -8361
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p35_Z5USRC  sky130_fd_pr__res_xhigh_po_0p35_Z5USRC_0
timestamp 1724926688
transform -1 0 25341 0 -1 -8361
box -699 -682 699 682
use sky130_fd_pr__res_xhigh_po_0p69_PWEJ5Z  sky130_fd_pr__res_xhigh_po_0p69_PWEJ5Z_0
timestamp 1724926688
transform 1 0 24557 0 1 -9834
box -1522 -708 1522 708
use sky130_fd_pr__pfet_01v8_lvt_6GTY34  XM1
timestamp 1724939774
transform 1 0 25356 0 1 -5820
box -855 -1098 855 1064
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2 ~/pdk/sky130A/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 5 1288
timestamp 1704896540
transform -1 0 33095 0 -1 -4445
box 0 0 1340 1340
<< labels >>
flabel metal2 19700 -6239 19796 -6064 0 FreeSans 160 0 0 0 Gcm1
port 3 nsew
flabel metal1 21001 -7152 21109 -7078 0 FreeSans 160 0 0 0 opout
port 8 nsew
flabel metal1 26176 -8411 26288 -8297 0 FreeSans 160 0 0 0 Vbgr
flabel metal1 20300 -9273 20400 -9211 0 FreeSans 160 0 0 0 Gcm2
port 4 nsew
flabel metal1 19841 -9319 19901 -9273 0 FreeSans 160 0 0 0 Sop
port 7 nsew
flabel metal1 22344 -4599 22547 -4401 0 FreeSans 160 0 0 0 Vbgr
port 9 nsew
flabel space 20000 -7806 20102 -7657 0 FreeSans 160 0 0 0 MINUS
port 6 nsew
flabel space 23298 -6830 23402 -6775 0 FreeSans 160 0 0 0 VSS
port 2 nsew
flabel metal3 20524 -4594 20654 -4534 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel space 19702 -7802 19804 -7654 0 FreeSans 160 0 0 0 PLUS
port 5 nsew
<< end >>
