** sch_path: /home/ttuser/tt08-bgr/xschem/PLSIM.sch
**.subckt PLSIM
V2 VSS GND 0
R1 Vbgr VSS 11G m=1
x1 VDD Vbgr VSS core_prel
R2 Vbgr_parax VSS 11G m=1
x2 VDD Vbgr_parax VSS core_prel_parax
V3 net1 VSS pwl 0 0 1u 0 4u VDD
E5 TEMPERAT VSS VOL=' temper '
.save v(temperat)
VDD net1 VDD 0
.save i(vdd)
.save v(vbgr)
.save v(vbgr_parax)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt




* this experimental option enables mos model bin
* selection based on W/NF instead of W
.options wnflag=1 XMU=0.49 METHOD=GEAR ITL4=100 CHGTOL=1e-15 TRTOL=1 RELTOL=0.0001 VNTOL=0.1u
.param ABSVAR=0.03
.param VCCGAUSS=agauss(1.8, 'ABSVAR', 1)
.param VDD=VCCGAUSS
*.param VDD=1.8
** variation marameters:
* .options savecurrents
.control
  setseed 12
  reset
  let run=1
  dowhile run <= 100
    if run > 1
      reset
      set appendwrite
    end
    * save all
    if run % 3 = 1
      set temp=-40
    end
    if run % 3 = 2
      set temp=27
    end
    if run % 3 = 0
      set temp=125
    end
    echo "Run=$&run, Temp=$temp"
    tran 0.2u 50u
    write plsim.raw
    let run = run + 1
  end
.endc


**** end user architecture code
**.ends

* expanding   symbol:  core_prel.sym # of pins=3
** sym_path: /home/ttuser/tt08-bgr/xschem/core_prel.sym
** sch_path: /home/ttuser/tt08-bgr/xschem/core_prel.sch
.subckt core_prel VDD Vbgr VSS
*.ipin VDD
*.ipin VSS
*.opin Vbgr
XQ1 VSS VSS MINUS sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ2 VSS VSS net1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=29
XM1 MINUS opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 PLUS opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vbgr opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 opout MINUS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Gcm1 PLUS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 opout Gcm1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 Sop Gcm2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 Gcm2 Gcm2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Gcm1 Gcm1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 Gcm2 opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR19 net1 PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=0.9 mult=1 m=1
XR3 VSS MINUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6 mult=1 m=1
XR4 VSS Vbgr VSS sky130_fd_pr__res_xhigh_po_0p69 L=12.6 mult=1 m=1
XM12 VSS Vbgr opout opout sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XR2 VSS PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6 mult=1 m=1
XM11 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR1 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p69 L=1.26 mult=1 m=1
XR5 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p69 L=1.26 mult=1 m=1
XR6 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
XR7 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
XM14 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 Gcm2 VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  core_prel_parax.sym # of pins=3
** sym_path: /home/ttuser/tt08-bgr/xschem/core_prel.sym
.include /home/ttuser/tt08-bgr/mag/core_prel.sim.spice
.GLOBAL GND
.end
