magic
tech sky130A
magscale 1 2
timestamp 1725004556
<< nwell >>
rect -1196 -973 1196 973
<< pmoslvt >>
rect -1000 554 1000 754
rect -1000 118 1000 318
rect -1000 -318 1000 -118
rect -1000 -754 1000 -554
<< pdiff >>
rect -1058 742 -1000 754
rect -1058 566 -1046 742
rect -1012 566 -1000 742
rect -1058 554 -1000 566
rect 1000 742 1058 754
rect 1000 566 1012 742
rect 1046 566 1058 742
rect 1000 554 1058 566
rect -1058 306 -1000 318
rect -1058 130 -1046 306
rect -1012 130 -1000 306
rect -1058 118 -1000 130
rect 1000 306 1058 318
rect 1000 130 1012 306
rect 1046 130 1058 306
rect 1000 118 1058 130
rect -1058 -130 -1000 -118
rect -1058 -306 -1046 -130
rect -1012 -306 -1000 -130
rect -1058 -318 -1000 -306
rect 1000 -130 1058 -118
rect 1000 -306 1012 -130
rect 1046 -306 1058 -130
rect 1000 -318 1058 -306
rect -1058 -566 -1000 -554
rect -1058 -742 -1046 -566
rect -1012 -742 -1000 -566
rect -1058 -754 -1000 -742
rect 1000 -566 1058 -554
rect 1000 -742 1012 -566
rect 1046 -742 1058 -566
rect 1000 -754 1058 -742
<< pdiffc >>
rect -1046 566 -1012 742
rect 1012 566 1046 742
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
rect -1046 -742 -1012 -566
rect 1012 -742 1046 -566
<< nsubdiff >>
rect -1160 903 1160 937
rect -1160 -903 -1126 903
rect 1126 841 1160 903
rect 1126 -903 1160 -841
rect -1160 -937 1160 -903
<< nsubdiffcont >>
rect 1126 -841 1160 841
<< poly >>
rect -1000 835 1000 851
rect -1000 801 -984 835
rect 984 801 1000 835
rect -1000 754 1000 801
rect -1000 507 1000 554
rect -1000 473 -984 507
rect 984 473 1000 507
rect -1000 457 1000 473
rect -1000 399 1000 415
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1000 318 1000 365
rect -1000 71 1000 118
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 21 1000 37
rect -1000 -37 1000 -21
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1000 -118 1000 -71
rect -1000 -365 1000 -318
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1000 -415 1000 -399
rect -1000 -473 1000 -457
rect -1000 -507 -984 -473
rect 984 -507 1000 -473
rect -1000 -554 1000 -507
rect -1000 -801 1000 -754
rect -1000 -835 -984 -801
rect 984 -835 1000 -801
rect -1000 -851 1000 -835
<< polycont >>
rect -984 801 984 835
rect -984 473 984 507
rect -984 365 984 399
rect -984 37 984 71
rect -984 -71 984 -37
rect -984 -399 984 -365
rect -984 -507 984 -473
rect -984 -835 984 -801
<< locali >>
rect 1126 841 1160 857
rect -1000 801 -984 835
rect 984 801 1000 835
rect -1046 742 -1012 758
rect -1046 550 -1012 566
rect 1012 742 1046 758
rect 1012 550 1046 566
rect -1000 473 -984 507
rect 984 473 1000 507
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1046 306 -1012 322
rect -1046 114 -1012 130
rect 1012 306 1046 322
rect 1012 114 1046 130
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1046 -130 -1012 -114
rect -1046 -322 -1012 -306
rect 1012 -130 1046 -114
rect 1012 -322 1046 -306
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1000 -507 -984 -473
rect 984 -507 1000 -473
rect -1046 -566 -1012 -550
rect -1046 -758 -1012 -742
rect 1012 -566 1046 -550
rect 1012 -758 1046 -742
rect -1000 -835 -984 -801
rect 984 -835 1000 -801
rect 1126 -857 1160 -841
<< viali >>
rect -492 801 492 835
rect -1046 566 -1012 742
rect 1012 566 1046 742
rect -492 473 492 507
rect -492 365 492 399
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -492 37 492 71
rect -492 -71 492 -37
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
rect -492 -399 492 -365
rect -492 -507 492 -473
rect -1046 -742 -1012 -566
rect 1012 -742 1046 -566
rect -492 -835 492 -801
<< metal1 >>
rect -504 835 504 841
rect -504 801 -492 835
rect 492 801 504 835
rect -504 795 504 801
rect -1052 742 -1006 754
rect -1052 566 -1046 742
rect -1012 566 -1006 742
rect -1052 554 -1006 566
rect 1006 742 1052 754
rect 1006 566 1012 742
rect 1046 566 1052 742
rect 1006 554 1052 566
rect -504 507 504 513
rect -504 473 -492 507
rect 492 473 504 507
rect -504 467 504 473
rect -504 399 504 405
rect -504 365 -492 399
rect 492 365 504 399
rect -504 359 504 365
rect -1052 306 -1006 318
rect -1052 130 -1046 306
rect -1012 130 -1006 306
rect -1052 118 -1006 130
rect 1006 306 1052 318
rect 1006 130 1012 306
rect 1046 130 1052 306
rect 1006 118 1052 130
rect -504 71 504 77
rect -504 37 -492 71
rect 492 37 504 71
rect -504 31 504 37
rect -504 -37 504 -31
rect -504 -71 -492 -37
rect 492 -71 504 -37
rect -504 -77 504 -71
rect -1052 -130 -1006 -118
rect -1052 -306 -1046 -130
rect -1012 -306 -1006 -130
rect -1052 -318 -1006 -306
rect 1006 -130 1052 -118
rect 1006 -306 1012 -130
rect 1046 -306 1052 -130
rect 1006 -318 1052 -306
rect -504 -365 504 -359
rect -504 -399 -492 -365
rect 492 -399 504 -365
rect -504 -405 504 -399
rect -504 -473 504 -467
rect -504 -507 -492 -473
rect 492 -507 504 -473
rect -504 -513 504 -507
rect -1052 -566 -1006 -554
rect -1052 -742 -1046 -566
rect -1012 -742 -1006 -566
rect -1052 -754 -1006 -742
rect 1006 -566 1052 -554
rect 1006 -742 1012 -566
rect 1046 -742 1052 -566
rect 1006 -754 1052 -742
rect -504 -801 504 -795
rect -504 -835 -492 -801
rect 492 -835 504 -801
rect -504 -841 504 -835
<< properties >>
string FIXED_BBOX -1143 -920 1143 920
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 10 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
