magic
tech sky130A
magscale 1 2
timestamp 1724543890
<< pwell >>
rect -201 -1217 201 1217
<< psubdiff >>
rect -165 1147 -69 1181
rect 69 1147 165 1181
rect -165 1085 -131 1147
rect 131 1085 165 1147
rect -165 -1147 -131 -1085
rect 131 -1147 165 -1085
rect -165 -1181 -69 -1147
rect 69 -1181 165 -1147
<< psubdiffcont >>
rect -69 1147 69 1181
rect -165 -1085 -131 1085
rect 131 -1085 165 1085
rect -69 -1181 69 -1147
<< xpolycontact >>
rect -35 619 35 1051
rect -35 -1051 35 -619
<< xpolyres >>
rect -35 -619 35 619
<< locali >>
rect -165 1147 -69 1181
rect 69 1147 165 1181
rect -165 1085 -131 1147
rect 131 1085 165 1147
rect -165 -1147 -131 -1085
rect 131 -1147 165 -1085
rect -165 -1181 -69 -1147
rect 69 -1181 165 -1147
<< viali >>
rect -19 636 19 1033
rect -19 -1033 19 -636
<< metal1 >>
rect -25 1033 25 1045
rect -25 636 -19 1033
rect 19 636 25 1033
rect -25 624 25 636
rect -25 -636 25 -624
rect -25 -1033 -19 -636
rect 19 -1033 25 -636
rect -25 -1045 25 -1033
<< properties >>
string FIXED_BBOX -148 -1164 148 1164
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 6.35 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 37.361k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
