magic
tech sky130A
magscale 1 2
timestamp 1724543890
<< pwell >>
rect -201 -675 201 675
<< psubdiff >>
rect -165 605 -69 639
rect 69 605 165 639
rect -165 543 -131 605
rect 131 543 165 605
rect -165 -605 -131 -543
rect 131 -605 165 -543
rect -165 -639 -69 -605
rect 69 -639 165 -605
<< psubdiffcont >>
rect -69 605 69 639
rect -165 -543 -131 543
rect 131 -543 165 543
rect -69 -639 69 -605
<< xpolycontact >>
rect -35 77 35 509
rect -35 -509 35 -77
<< xpolyres >>
rect -35 -77 35 77
<< locali >>
rect -165 605 -69 639
rect 69 605 165 639
rect -165 543 -131 605
rect 131 543 165 605
rect -165 -605 -131 -543
rect 131 -605 165 -543
rect -165 -639 -69 -605
rect 69 -639 165 -605
<< viali >>
rect -19 94 19 491
rect -19 -491 19 -94
<< metal1 >>
rect -25 491 25 503
rect -25 94 -19 491
rect 19 94 25 491
rect -25 82 25 94
rect -25 -94 25 -82
rect -25 -491 -19 -94
rect 19 -491 25 -94
rect -25 -503 25 -491
<< properties >>
string FIXED_BBOX -148 -622 148 622
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.93 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 6.389k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
