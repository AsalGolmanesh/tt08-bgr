** sch_path: /home/ttuser/tt08-bgr/xschem/BGRwOpampRes.sch
**.subckt BGRwOpampRes
XQ1 VSS VSS MINUS sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ2 VSS VSS net8 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=29
XM1 net1 vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vbgr vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V2 VSS GND 0
Vmeas net1 MINUS 0
.save i(vmeas)
Vmeas1 net2 PLUS 0
.save i(vmeas1)
.save v(vdd)
.save v(net1)
.save v(vdd)
.save v(net2)
.save v(vdd)
.save v(vbgr)
XM4 vp MINUS net3 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net5 PLUS net3 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 vp net5 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.save v(vp)
.save v(net3)
.save v(net5)
.save v(net3)
XM10 net6 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net5 net5 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.save v(vdd)
.save v(net5)
.save v(vdd)
.save v(vp)
.save v(net6)
.save v(vss)
.save v(net4)
.save v(vss)
Vmeas3 net3 net6 0
.save i(vmeas3)
XM8 net7 vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas2 net7 net4 0
.save i(vmeas2)
.save v(vdd)
.save v(net7)
XM11 VSS Vbgr vp vp sky130_fd_pr__pfet_01v8_lvt L=35 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V3 net9 VSS pwl 0 0 1u 0 4u VDD
E5 TEMPERAT VSS VOL=' temper '
.save v(temperat)
VDD net9 VDD 0
.save i(vdd)
.save v(minus)
.save v(plus)
XR19 net8 PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=0.93 mult=1 m=1
XR2 VSS PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6.35 mult=1 m=1
XR3 VSS MINUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6.35 mult=1 m=1
XR1 VSS Vbgr VSS sky130_fd_pr__res_xhigh_po_1p41 L=26.57 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt




* this experimental option enables mos model bin
* selection based on W/NF instead of W
* .options wnflag=1 XMU=0.49 METHOD=GEAR ITL4=100 CHGTOL=1e-15 TRTOL=1 RELTOL=0.0001 VNTOL=0.1u
.param ABSVAR=0.03
.param VCCGAUSS=agauss(1.8, 'ABSVAR', 1)
.param VDD=VCCGAUSS
*.param VDD=1.8
** variation marameters:
* .options savecurrents
.control
  setseed 12
  reset
  let run=1
  dowhile run <= 100
    if run > 1
      reset
      set appendwrite
    end
    * save all
    if run % 3 = 1
      set temp=-40
    end
    if run % 3 = 2
      set temp=27
    end
    if run % 3 = 0
      set temp=125
    end
    echo "Run=$&run, Temp=$temp"
    tran 0.2u 50u
    write asal_tb_bandgap_r.raw
    let run = run + 1
  end
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
